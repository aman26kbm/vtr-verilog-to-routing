`timescale 1ns/1ns
`define DWIDTH 16
`define AWIDTH 7
`define MEM_SIZE 128
`define BB_MAT_MUL_SIZE 4


module matrix_multiplication(
  clk,
  reset,
  enable_writing_to_mem,
  enable_reading_from_mem,
  data_pi,
  addr_pi,
  we_a,
  we_b,
  we_c,
  data_from_out_mat,
  start_mat_mul,
  done_mat_mul
);

  input clk;
  input reset;
  input enable_writing_to_mem;
  input enable_reading_from_mem;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_pi;
  input [`AWIDTH-1:0] addr_pi;
  input we_a;
  input we_b;
  input we_c;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat;
  input start_mat_mul;
  output done_mat_mul;



  reg enable_writing_to_mem_reg;
  reg [`AWIDTH-1:0] addr_pi_reg;
  always @(posedge clk) begin
    if (reset) begin
      enable_writing_to_mem_reg <= 0;
      addr_pi_reg <= 0;
    end else begin
      enable_writing_to_mem_reg <= enable_writing_to_mem;
      addr_pi_reg <= addr_pi;
    end
  end
/////////////////////////////////////////////////
// BRAMs to store matrix A
/////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_0;
  wire [`AWIDTH-1:0] a_addr_0_0;
  wire [`AWIDTH-1:0] a_addr_muxed_0_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_0_0_reg;
  reg  [`AWIDTH-1:0] a_addr_0_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_0_0_reg <= 0;
      a_addr_muxed_0_0_reg <= 0;
    end else begin
      a_addr_0_0_reg <= a_addr_0_0;
      a_addr_muxed_0_0_reg <= a_addr_muxed_0_0;
    end
  end
  assign a_addr_muxed_0_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_0_0_reg;

  // BRAM matrix A 0_0
  ram matrix_A_0_0 (
    .addr0(a_addr_muxed_0_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_0_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_0;
  wire [`AWIDTH-1:0] a_addr_1_0;
  wire [`AWIDTH-1:0] a_addr_muxed_1_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_1_0_reg;
  reg  [`AWIDTH-1:0] a_addr_1_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_1_0_reg <= 0;
      a_addr_muxed_1_0_reg <= 0;
    end else begin
      a_addr_1_0_reg <= a_addr_1_0;
      a_addr_muxed_1_0_reg <= a_addr_muxed_1_0;
    end
  end
  assign a_addr_muxed_1_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_1_0_reg;

  // BRAM matrix A 1_0
  ram matrix_A_1_0 (
    .addr0(a_addr_muxed_1_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_1_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_0;
  wire [`AWIDTH-1:0] a_addr_2_0;
  wire [`AWIDTH-1:0] a_addr_muxed_2_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_2_0_reg;
  reg  [`AWIDTH-1:0] a_addr_2_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_2_0_reg <= 0;
      a_addr_muxed_2_0_reg <= 0;
    end else begin
      a_addr_2_0_reg <= a_addr_2_0;
      a_addr_muxed_2_0_reg <= a_addr_muxed_2_0;
    end
  end
  assign a_addr_muxed_2_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_2_0_reg;

  // BRAM matrix A 2_0
  ram matrix_A_2_0 (
    .addr0(a_addr_muxed_2_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_2_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_0;
  wire [`AWIDTH-1:0] a_addr_3_0;
  wire [`AWIDTH-1:0] a_addr_muxed_3_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_3_0_reg;
  reg  [`AWIDTH-1:0] a_addr_3_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_3_0_reg <= 0;
      a_addr_muxed_3_0_reg <= 0;
    end else begin
      a_addr_3_0_reg <= a_addr_3_0;
      a_addr_muxed_3_0_reg <= a_addr_muxed_3_0;
    end
  end
  assign a_addr_muxed_3_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_3_0_reg;

  // BRAM matrix A 3_0
  ram matrix_A_3_0 (
    .addr0(a_addr_muxed_3_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_3_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_0;
  wire [`AWIDTH-1:0] a_addr_4_0;
  wire [`AWIDTH-1:0] a_addr_muxed_4_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_4_0_reg;
  reg  [`AWIDTH-1:0] a_addr_4_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_4_0_reg <= 0;
      a_addr_muxed_4_0_reg <= 0;
    end else begin
      a_addr_4_0_reg <= a_addr_4_0;
      a_addr_muxed_4_0_reg <= a_addr_muxed_4_0;
    end
  end
  assign a_addr_muxed_4_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_4_0_reg;

  // BRAM matrix A 4_0
  ram matrix_A_4_0 (
    .addr0(a_addr_muxed_4_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_4_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_0;
  wire [`AWIDTH-1:0] a_addr_5_0;
  wire [`AWIDTH-1:0] a_addr_muxed_5_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_5_0_reg;
  reg  [`AWIDTH-1:0] a_addr_5_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_5_0_reg <= 0;
      a_addr_muxed_5_0_reg <= 0;
    end else begin
      a_addr_5_0_reg <= a_addr_5_0;
      a_addr_muxed_5_0_reg <= a_addr_muxed_5_0;
    end
  end
  assign a_addr_muxed_5_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_5_0_reg;

  // BRAM matrix A 5_0
  ram matrix_A_5_0 (
    .addr0(a_addr_muxed_5_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_5_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_0;
  wire [`AWIDTH-1:0] a_addr_6_0;
  wire [`AWIDTH-1:0] a_addr_muxed_6_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_6_0_reg;
  reg  [`AWIDTH-1:0] a_addr_6_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_6_0_reg <= 0;
      a_addr_muxed_6_0_reg <= 0;
    end else begin
      a_addr_6_0_reg <= a_addr_6_0;
      a_addr_muxed_6_0_reg <= a_addr_muxed_6_0;
    end
  end
  assign a_addr_muxed_6_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_6_0_reg;

  // BRAM matrix A 6_0
  ram matrix_A_6_0 (
    .addr0(a_addr_muxed_6_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_6_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_0;
  wire [`AWIDTH-1:0] a_addr_7_0;
  wire [`AWIDTH-1:0] a_addr_muxed_7_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_7_0_reg;
  reg  [`AWIDTH-1:0] a_addr_7_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_7_0_reg <= 0;
      a_addr_muxed_7_0_reg <= 0;
    end else begin
      a_addr_7_0_reg <= a_addr_7_0;
      a_addr_muxed_7_0_reg <= a_addr_muxed_7_0;
    end
  end
  assign a_addr_muxed_7_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_7_0_reg;

  // BRAM matrix A 7_0
  ram matrix_A_7_0 (
    .addr0(a_addr_muxed_7_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_7_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_0;
  wire [`AWIDTH-1:0] a_addr_8_0;
  wire [`AWIDTH-1:0] a_addr_muxed_8_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_8_0_reg;
  reg  [`AWIDTH-1:0] a_addr_8_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_8_0_reg <= 0;
      a_addr_muxed_8_0_reg <= 0;
    end else begin
      a_addr_8_0_reg <= a_addr_8_0;
      a_addr_muxed_8_0_reg <= a_addr_muxed_8_0;
    end
  end
  assign a_addr_muxed_8_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_8_0_reg;

  // BRAM matrix A 8_0
  ram matrix_A_8_0 (
    .addr0(a_addr_muxed_8_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_8_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_0;
  wire [`AWIDTH-1:0] a_addr_9_0;
  wire [`AWIDTH-1:0] a_addr_muxed_9_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_9_0_reg;
  reg  [`AWIDTH-1:0] a_addr_9_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_9_0_reg <= 0;
      a_addr_muxed_9_0_reg <= 0;
    end else begin
      a_addr_9_0_reg <= a_addr_9_0;
      a_addr_muxed_9_0_reg <= a_addr_muxed_9_0;
    end
  end
  assign a_addr_muxed_9_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_9_0_reg;

  // BRAM matrix A 9_0
  ram matrix_A_9_0 (
    .addr0(a_addr_muxed_9_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_9_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_0;
  wire [`AWIDTH-1:0] a_addr_10_0;
  wire [`AWIDTH-1:0] a_addr_muxed_10_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_10_0_reg;
  reg  [`AWIDTH-1:0] a_addr_10_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_10_0_reg <= 0;
      a_addr_muxed_10_0_reg <= 0;
    end else begin
      a_addr_10_0_reg <= a_addr_10_0;
      a_addr_muxed_10_0_reg <= a_addr_muxed_10_0;
    end
  end
  assign a_addr_muxed_10_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_10_0_reg;

  // BRAM matrix A 10_0
  ram matrix_A_10_0 (
    .addr0(a_addr_muxed_10_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_10_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_0;
  wire [`AWIDTH-1:0] a_addr_11_0;
  wire [`AWIDTH-1:0] a_addr_muxed_11_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_11_0_reg;
  reg  [`AWIDTH-1:0] a_addr_11_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_11_0_reg <= 0;
      a_addr_muxed_11_0_reg <= 0;
    end else begin
      a_addr_11_0_reg <= a_addr_11_0;
      a_addr_muxed_11_0_reg <= a_addr_muxed_11_0;
    end
  end
  assign a_addr_muxed_11_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_11_0_reg;

  // BRAM matrix A 11_0
  ram matrix_A_11_0 (
    .addr0(a_addr_muxed_11_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_11_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_0;
  wire [`AWIDTH-1:0] a_addr_12_0;
  wire [`AWIDTH-1:0] a_addr_muxed_12_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_12_0_reg;
  reg  [`AWIDTH-1:0] a_addr_12_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_12_0_reg <= 0;
      a_addr_muxed_12_0_reg <= 0;
    end else begin
      a_addr_12_0_reg <= a_addr_12_0;
      a_addr_muxed_12_0_reg <= a_addr_muxed_12_0;
    end
  end
  assign a_addr_muxed_12_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_12_0_reg;

  // BRAM matrix A 12_0
  ram matrix_A_12_0 (
    .addr0(a_addr_muxed_12_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_12_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_0;
  wire [`AWIDTH-1:0] a_addr_13_0;
  wire [`AWIDTH-1:0] a_addr_muxed_13_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_13_0_reg;
  reg  [`AWIDTH-1:0] a_addr_13_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_13_0_reg <= 0;
      a_addr_muxed_13_0_reg <= 0;
    end else begin
      a_addr_13_0_reg <= a_addr_13_0;
      a_addr_muxed_13_0_reg <= a_addr_muxed_13_0;
    end
  end
  assign a_addr_muxed_13_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_13_0_reg;

  // BRAM matrix A 13_0
  ram matrix_A_13_0 (
    .addr0(a_addr_muxed_13_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_13_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_0;
  wire [`AWIDTH-1:0] a_addr_14_0;
  wire [`AWIDTH-1:0] a_addr_muxed_14_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_14_0_reg;
  reg  [`AWIDTH-1:0] a_addr_14_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_14_0_reg <= 0;
      a_addr_muxed_14_0_reg <= 0;
    end else begin
      a_addr_14_0_reg <= a_addr_14_0;
      a_addr_muxed_14_0_reg <= a_addr_muxed_14_0;
    end
  end
  assign a_addr_muxed_14_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_14_0_reg;

  // BRAM matrix A 14_0
  ram matrix_A_14_0 (
    .addr0(a_addr_muxed_14_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_14_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_0;
  wire [`AWIDTH-1:0] a_addr_15_0;
  wire [`AWIDTH-1:0] a_addr_muxed_15_0;

  reg  [`AWIDTH-1:0] a_addr_muxed_15_0_reg;
  reg  [`AWIDTH-1:0] a_addr_15_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      a_addr_15_0_reg <= 0;
      a_addr_muxed_15_0_reg <= 0;
    end else begin
      a_addr_15_0_reg <= a_addr_15_0;
      a_addr_muxed_15_0_reg <= a_addr_muxed_15_0;
    end
  end
  assign a_addr_muxed_15_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : a_addr_15_0_reg;

  // BRAM matrix A 15_0
  ram matrix_A_15_0 (
    .addr0(a_addr_muxed_15_0_reg),
    .d0(data_pi),
    .we0(we_a),
    .q0(a_data_15_0),
    .clk(clk));

/////////////////////////////////////////////////
// BRAMs to store matrix B
/////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_0;
  wire [`AWIDTH-1:0] b_addr_0_0;
  wire [`AWIDTH-1:0] b_addr_muxed_0_0;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_0_reg;
  reg  [`AWIDTH-1:0] b_addr_0_0_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_0_reg <= 0;
      b_addr_muxed_0_0_reg <= 0;
    end else begin
      b_addr_0_0_reg <= b_addr_0_0;
      b_addr_muxed_0_0_reg <= b_addr_muxed_0_0;
    end
  end
  assign b_addr_muxed_0_0 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_0_reg;

  // BRAM matrix B 0_0
  ram matrix_B_0_0 (
    .addr0(b_addr_muxed_0_0_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_0),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_1;
  wire [`AWIDTH-1:0] b_addr_0_1;
  wire [`AWIDTH-1:0] b_addr_muxed_0_1;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_1_reg;
  reg  [`AWIDTH-1:0] b_addr_0_1_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_1_reg <= 0;
      b_addr_muxed_0_1_reg <= 0;
    end else begin
      b_addr_0_1_reg <= b_addr_0_1;
      b_addr_muxed_0_1_reg <= b_addr_muxed_0_1;
    end
  end
  assign b_addr_muxed_0_1 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_1_reg;

  // BRAM matrix B 0_1
  ram matrix_B_0_1 (
    .addr0(b_addr_muxed_0_1_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_1),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_2;
  wire [`AWIDTH-1:0] b_addr_0_2;
  wire [`AWIDTH-1:0] b_addr_muxed_0_2;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_2_reg;
  reg  [`AWIDTH-1:0] b_addr_0_2_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_2_reg <= 0;
      b_addr_muxed_0_2_reg <= 0;
    end else begin
      b_addr_0_2_reg <= b_addr_0_2;
      b_addr_muxed_0_2_reg <= b_addr_muxed_0_2;
    end
  end
  assign b_addr_muxed_0_2 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_2_reg;

  // BRAM matrix B 0_2
  ram matrix_B_0_2 (
    .addr0(b_addr_muxed_0_2_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_2),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_3;
  wire [`AWIDTH-1:0] b_addr_0_3;
  wire [`AWIDTH-1:0] b_addr_muxed_0_3;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_3_reg;
  reg  [`AWIDTH-1:0] b_addr_0_3_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_3_reg <= 0;
      b_addr_muxed_0_3_reg <= 0;
    end else begin
      b_addr_0_3_reg <= b_addr_0_3;
      b_addr_muxed_0_3_reg <= b_addr_muxed_0_3;
    end
  end
  assign b_addr_muxed_0_3 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_3_reg;

  // BRAM matrix B 0_3
  ram matrix_B_0_3 (
    .addr0(b_addr_muxed_0_3_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_3),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_4;
  wire [`AWIDTH-1:0] b_addr_0_4;
  wire [`AWIDTH-1:0] b_addr_muxed_0_4;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_4_reg;
  reg  [`AWIDTH-1:0] b_addr_0_4_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_4_reg <= 0;
      b_addr_muxed_0_4_reg <= 0;
    end else begin
      b_addr_0_4_reg <= b_addr_0_4;
      b_addr_muxed_0_4_reg <= b_addr_muxed_0_4;
    end
  end
  assign b_addr_muxed_0_4 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_4_reg;

  // BRAM matrix B 0_4
  ram matrix_B_0_4 (
    .addr0(b_addr_muxed_0_4_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_4),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_5;
  wire [`AWIDTH-1:0] b_addr_0_5;
  wire [`AWIDTH-1:0] b_addr_muxed_0_5;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_5_reg;
  reg  [`AWIDTH-1:0] b_addr_0_5_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_5_reg <= 0;
      b_addr_muxed_0_5_reg <= 0;
    end else begin
      b_addr_0_5_reg <= b_addr_0_5;
      b_addr_muxed_0_5_reg <= b_addr_muxed_0_5;
    end
  end
  assign b_addr_muxed_0_5 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_5_reg;

  // BRAM matrix B 0_5
  ram matrix_B_0_5 (
    .addr0(b_addr_muxed_0_5_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_5),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_6;
  wire [`AWIDTH-1:0] b_addr_0_6;
  wire [`AWIDTH-1:0] b_addr_muxed_0_6;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_6_reg;
  reg  [`AWIDTH-1:0] b_addr_0_6_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_6_reg <= 0;
      b_addr_muxed_0_6_reg <= 0;
    end else begin
      b_addr_0_6_reg <= b_addr_0_6;
      b_addr_muxed_0_6_reg <= b_addr_muxed_0_6;
    end
  end
  assign b_addr_muxed_0_6 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_6_reg;

  // BRAM matrix B 0_6
  ram matrix_B_0_6 (
    .addr0(b_addr_muxed_0_6_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_6),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_7;
  wire [`AWIDTH-1:0] b_addr_0_7;
  wire [`AWIDTH-1:0] b_addr_muxed_0_7;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_7_reg;
  reg  [`AWIDTH-1:0] b_addr_0_7_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_7_reg <= 0;
      b_addr_muxed_0_7_reg <= 0;
    end else begin
      b_addr_0_7_reg <= b_addr_0_7;
      b_addr_muxed_0_7_reg <= b_addr_muxed_0_7;
    end
  end
  assign b_addr_muxed_0_7 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_7_reg;

  // BRAM matrix B 0_7
  ram matrix_B_0_7 (
    .addr0(b_addr_muxed_0_7_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_7),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_8;
  wire [`AWIDTH-1:0] b_addr_0_8;
  wire [`AWIDTH-1:0] b_addr_muxed_0_8;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_8_reg;
  reg  [`AWIDTH-1:0] b_addr_0_8_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_8_reg <= 0;
      b_addr_muxed_0_8_reg <= 0;
    end else begin
      b_addr_0_8_reg <= b_addr_0_8;
      b_addr_muxed_0_8_reg <= b_addr_muxed_0_8;
    end
  end
  assign b_addr_muxed_0_8 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_8_reg;

  // BRAM matrix B 0_8
  ram matrix_B_0_8 (
    .addr0(b_addr_muxed_0_8_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_8),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_9;
  wire [`AWIDTH-1:0] b_addr_0_9;
  wire [`AWIDTH-1:0] b_addr_muxed_0_9;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_9_reg;
  reg  [`AWIDTH-1:0] b_addr_0_9_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_9_reg <= 0;
      b_addr_muxed_0_9_reg <= 0;
    end else begin
      b_addr_0_9_reg <= b_addr_0_9;
      b_addr_muxed_0_9_reg <= b_addr_muxed_0_9;
    end
  end
  assign b_addr_muxed_0_9 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_9_reg;

  // BRAM matrix B 0_9
  ram matrix_B_0_9 (
    .addr0(b_addr_muxed_0_9_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_9),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_10;
  wire [`AWIDTH-1:0] b_addr_0_10;
  wire [`AWIDTH-1:0] b_addr_muxed_0_10;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_10_reg;
  reg  [`AWIDTH-1:0] b_addr_0_10_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_10_reg <= 0;
      b_addr_muxed_0_10_reg <= 0;
    end else begin
      b_addr_0_10_reg <= b_addr_0_10;
      b_addr_muxed_0_10_reg <= b_addr_muxed_0_10;
    end
  end
  assign b_addr_muxed_0_10 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_10_reg;

  // BRAM matrix B 0_10
  ram matrix_B_0_10 (
    .addr0(b_addr_muxed_0_10_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_10),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_11;
  wire [`AWIDTH-1:0] b_addr_0_11;
  wire [`AWIDTH-1:0] b_addr_muxed_0_11;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_11_reg;
  reg  [`AWIDTH-1:0] b_addr_0_11_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_11_reg <= 0;
      b_addr_muxed_0_11_reg <= 0;
    end else begin
      b_addr_0_11_reg <= b_addr_0_11;
      b_addr_muxed_0_11_reg <= b_addr_muxed_0_11;
    end
  end
  assign b_addr_muxed_0_11 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_11_reg;

  // BRAM matrix B 0_11
  ram matrix_B_0_11 (
    .addr0(b_addr_muxed_0_11_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_11),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_12;
  wire [`AWIDTH-1:0] b_addr_0_12;
  wire [`AWIDTH-1:0] b_addr_muxed_0_12;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_12_reg;
  reg  [`AWIDTH-1:0] b_addr_0_12_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_12_reg <= 0;
      b_addr_muxed_0_12_reg <= 0;
    end else begin
      b_addr_0_12_reg <= b_addr_0_12;
      b_addr_muxed_0_12_reg <= b_addr_muxed_0_12;
    end
  end
  assign b_addr_muxed_0_12 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_12_reg;

  // BRAM matrix B 0_12
  ram matrix_B_0_12 (
    .addr0(b_addr_muxed_0_12_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_12),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_13;
  wire [`AWIDTH-1:0] b_addr_0_13;
  wire [`AWIDTH-1:0] b_addr_muxed_0_13;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_13_reg;
  reg  [`AWIDTH-1:0] b_addr_0_13_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_13_reg <= 0;
      b_addr_muxed_0_13_reg <= 0;
    end else begin
      b_addr_0_13_reg <= b_addr_0_13;
      b_addr_muxed_0_13_reg <= b_addr_muxed_0_13;
    end
  end
  assign b_addr_muxed_0_13 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_13_reg;

  // BRAM matrix B 0_13
  ram matrix_B_0_13 (
    .addr0(b_addr_muxed_0_13_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_13),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_14;
  wire [`AWIDTH-1:0] b_addr_0_14;
  wire [`AWIDTH-1:0] b_addr_muxed_0_14;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_14_reg;
  reg  [`AWIDTH-1:0] b_addr_0_14_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_14_reg <= 0;
      b_addr_muxed_0_14_reg <= 0;
    end else begin
      b_addr_0_14_reg <= b_addr_0_14;
      b_addr_muxed_0_14_reg <= b_addr_muxed_0_14;
    end
  end
  assign b_addr_muxed_0_14 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_14_reg;

  // BRAM matrix B 0_14
  ram matrix_B_0_14 (
    .addr0(b_addr_muxed_0_14_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_14),
    .clk(clk));

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_15;
  wire [`AWIDTH-1:0] b_addr_0_15;
  wire [`AWIDTH-1:0] b_addr_muxed_0_15;

  reg  [`AWIDTH-1:0] b_addr_muxed_0_15_reg;
  reg  [`AWIDTH-1:0] b_addr_0_15_reg;
  always @(posedge clk) begin
    if(reset) begin
      b_addr_0_15_reg <= 0;
      b_addr_muxed_0_15_reg <= 0;
    end else begin
      b_addr_0_15_reg <= b_addr_0_15;
      b_addr_muxed_0_15_reg <= b_addr_muxed_0_15;
    end
  end
  assign b_addr_muxed_0_15 = (enable_writing_to_mem_reg) ? addr_pi_reg : b_addr_0_15_reg;

  // BRAM matrix B 0_15
  ram matrix_B_0_15 (
    .addr0(b_addr_muxed_0_15_reg),
    .d0(data_pi),
    .we0(we_b),
    .q0(b_data_0_15),
    .clk(clk));

/////////////////////////////////////////////////
// BRAMs to store matrix C
/////////////////////////////////////////////////

  wire [`AWIDTH-1:0] c_addr_0_0;
  wire [`AWIDTH-1:0] c_addr_0_1;
  wire [`AWIDTH-1:0] c_addr_0_2;
  wire [`AWIDTH-1:0] c_addr_0_3;
  wire [`AWIDTH-1:0] c_addr_0_4;
  wire [`AWIDTH-1:0] c_addr_0_5;
  wire [`AWIDTH-1:0] c_addr_0_6;
  wire [`AWIDTH-1:0] c_addr_0_7;
  wire [`AWIDTH-1:0] c_addr_0_8;
  wire [`AWIDTH-1:0] c_addr_0_9;
  wire [`AWIDTH-1:0] c_addr_0_10;
  wire [`AWIDTH-1:0] c_addr_0_11;
  wire [`AWIDTH-1:0] c_addr_0_12;
  wire [`AWIDTH-1:0] c_addr_0_13;
  wire [`AWIDTH-1:0] c_addr_0_14;
  wire [`AWIDTH-1:0] c_addr_0_15;
  wire [`AWIDTH-1:0] c_addr_1_0;
  wire [`AWIDTH-1:0] c_addr_1_1;
  wire [`AWIDTH-1:0] c_addr_1_2;
  wire [`AWIDTH-1:0] c_addr_1_3;
  wire [`AWIDTH-1:0] c_addr_1_4;
  wire [`AWIDTH-1:0] c_addr_1_5;
  wire [`AWIDTH-1:0] c_addr_1_6;
  wire [`AWIDTH-1:0] c_addr_1_7;
  wire [`AWIDTH-1:0] c_addr_1_8;
  wire [`AWIDTH-1:0] c_addr_1_9;
  wire [`AWIDTH-1:0] c_addr_1_10;
  wire [`AWIDTH-1:0] c_addr_1_11;
  wire [`AWIDTH-1:0] c_addr_1_12;
  wire [`AWIDTH-1:0] c_addr_1_13;
  wire [`AWIDTH-1:0] c_addr_1_14;
  wire [`AWIDTH-1:0] c_addr_1_15;
  wire [`AWIDTH-1:0] c_addr_2_0;
  wire [`AWIDTH-1:0] c_addr_2_1;
  wire [`AWIDTH-1:0] c_addr_2_2;
  wire [`AWIDTH-1:0] c_addr_2_3;
  wire [`AWIDTH-1:0] c_addr_2_4;
  wire [`AWIDTH-1:0] c_addr_2_5;
  wire [`AWIDTH-1:0] c_addr_2_6;
  wire [`AWIDTH-1:0] c_addr_2_7;
  wire [`AWIDTH-1:0] c_addr_2_8;
  wire [`AWIDTH-1:0] c_addr_2_9;
  wire [`AWIDTH-1:0] c_addr_2_10;
  wire [`AWIDTH-1:0] c_addr_2_11;
  wire [`AWIDTH-1:0] c_addr_2_12;
  wire [`AWIDTH-1:0] c_addr_2_13;
  wire [`AWIDTH-1:0] c_addr_2_14;
  wire [`AWIDTH-1:0] c_addr_2_15;
  wire [`AWIDTH-1:0] c_addr_3_0;
  wire [`AWIDTH-1:0] c_addr_3_1;
  wire [`AWIDTH-1:0] c_addr_3_2;
  wire [`AWIDTH-1:0] c_addr_3_3;
  wire [`AWIDTH-1:0] c_addr_3_4;
  wire [`AWIDTH-1:0] c_addr_3_5;
  wire [`AWIDTH-1:0] c_addr_3_6;
  wire [`AWIDTH-1:0] c_addr_3_7;
  wire [`AWIDTH-1:0] c_addr_3_8;
  wire [`AWIDTH-1:0] c_addr_3_9;
  wire [`AWIDTH-1:0] c_addr_3_10;
  wire [`AWIDTH-1:0] c_addr_3_11;
  wire [`AWIDTH-1:0] c_addr_3_12;
  wire [`AWIDTH-1:0] c_addr_3_13;
  wire [`AWIDTH-1:0] c_addr_3_14;
  wire [`AWIDTH-1:0] c_addr_3_15;
  wire [`AWIDTH-1:0] c_addr_4_0;
  wire [`AWIDTH-1:0] c_addr_4_1;
  wire [`AWIDTH-1:0] c_addr_4_2;
  wire [`AWIDTH-1:0] c_addr_4_3;
  wire [`AWIDTH-1:0] c_addr_4_4;
  wire [`AWIDTH-1:0] c_addr_4_5;
  wire [`AWIDTH-1:0] c_addr_4_6;
  wire [`AWIDTH-1:0] c_addr_4_7;
  wire [`AWIDTH-1:0] c_addr_4_8;
  wire [`AWIDTH-1:0] c_addr_4_9;
  wire [`AWIDTH-1:0] c_addr_4_10;
  wire [`AWIDTH-1:0] c_addr_4_11;
  wire [`AWIDTH-1:0] c_addr_4_12;
  wire [`AWIDTH-1:0] c_addr_4_13;
  wire [`AWIDTH-1:0] c_addr_4_14;
  wire [`AWIDTH-1:0] c_addr_4_15;
  wire [`AWIDTH-1:0] c_addr_5_0;
  wire [`AWIDTH-1:0] c_addr_5_1;
  wire [`AWIDTH-1:0] c_addr_5_2;
  wire [`AWIDTH-1:0] c_addr_5_3;
  wire [`AWIDTH-1:0] c_addr_5_4;
  wire [`AWIDTH-1:0] c_addr_5_5;
  wire [`AWIDTH-1:0] c_addr_5_6;
  wire [`AWIDTH-1:0] c_addr_5_7;
  wire [`AWIDTH-1:0] c_addr_5_8;
  wire [`AWIDTH-1:0] c_addr_5_9;
  wire [`AWIDTH-1:0] c_addr_5_10;
  wire [`AWIDTH-1:0] c_addr_5_11;
  wire [`AWIDTH-1:0] c_addr_5_12;
  wire [`AWIDTH-1:0] c_addr_5_13;
  wire [`AWIDTH-1:0] c_addr_5_14;
  wire [`AWIDTH-1:0] c_addr_5_15;
  wire [`AWIDTH-1:0] c_addr_6_0;
  wire [`AWIDTH-1:0] c_addr_6_1;
  wire [`AWIDTH-1:0] c_addr_6_2;
  wire [`AWIDTH-1:0] c_addr_6_3;
  wire [`AWIDTH-1:0] c_addr_6_4;
  wire [`AWIDTH-1:0] c_addr_6_5;
  wire [`AWIDTH-1:0] c_addr_6_6;
  wire [`AWIDTH-1:0] c_addr_6_7;
  wire [`AWIDTH-1:0] c_addr_6_8;
  wire [`AWIDTH-1:0] c_addr_6_9;
  wire [`AWIDTH-1:0] c_addr_6_10;
  wire [`AWIDTH-1:0] c_addr_6_11;
  wire [`AWIDTH-1:0] c_addr_6_12;
  wire [`AWIDTH-1:0] c_addr_6_13;
  wire [`AWIDTH-1:0] c_addr_6_14;
  wire [`AWIDTH-1:0] c_addr_6_15;
  wire [`AWIDTH-1:0] c_addr_7_0;
  wire [`AWIDTH-1:0] c_addr_7_1;
  wire [`AWIDTH-1:0] c_addr_7_2;
  wire [`AWIDTH-1:0] c_addr_7_3;
  wire [`AWIDTH-1:0] c_addr_7_4;
  wire [`AWIDTH-1:0] c_addr_7_5;
  wire [`AWIDTH-1:0] c_addr_7_6;
  wire [`AWIDTH-1:0] c_addr_7_7;
  wire [`AWIDTH-1:0] c_addr_7_8;
  wire [`AWIDTH-1:0] c_addr_7_9;
  wire [`AWIDTH-1:0] c_addr_7_10;
  wire [`AWIDTH-1:0] c_addr_7_11;
  wire [`AWIDTH-1:0] c_addr_7_12;
  wire [`AWIDTH-1:0] c_addr_7_13;
  wire [`AWIDTH-1:0] c_addr_7_14;
  wire [`AWIDTH-1:0] c_addr_7_15;
  wire [`AWIDTH-1:0] c_addr_8_0;
  wire [`AWIDTH-1:0] c_addr_8_1;
  wire [`AWIDTH-1:0] c_addr_8_2;
  wire [`AWIDTH-1:0] c_addr_8_3;
  wire [`AWIDTH-1:0] c_addr_8_4;
  wire [`AWIDTH-1:0] c_addr_8_5;
  wire [`AWIDTH-1:0] c_addr_8_6;
  wire [`AWIDTH-1:0] c_addr_8_7;
  wire [`AWIDTH-1:0] c_addr_8_8;
  wire [`AWIDTH-1:0] c_addr_8_9;
  wire [`AWIDTH-1:0] c_addr_8_10;
  wire [`AWIDTH-1:0] c_addr_8_11;
  wire [`AWIDTH-1:0] c_addr_8_12;
  wire [`AWIDTH-1:0] c_addr_8_13;
  wire [`AWIDTH-1:0] c_addr_8_14;
  wire [`AWIDTH-1:0] c_addr_8_15;
  wire [`AWIDTH-1:0] c_addr_9_0;
  wire [`AWIDTH-1:0] c_addr_9_1;
  wire [`AWIDTH-1:0] c_addr_9_2;
  wire [`AWIDTH-1:0] c_addr_9_3;
  wire [`AWIDTH-1:0] c_addr_9_4;
  wire [`AWIDTH-1:0] c_addr_9_5;
  wire [`AWIDTH-1:0] c_addr_9_6;
  wire [`AWIDTH-1:0] c_addr_9_7;
  wire [`AWIDTH-1:0] c_addr_9_8;
  wire [`AWIDTH-1:0] c_addr_9_9;
  wire [`AWIDTH-1:0] c_addr_9_10;
  wire [`AWIDTH-1:0] c_addr_9_11;
  wire [`AWIDTH-1:0] c_addr_9_12;
  wire [`AWIDTH-1:0] c_addr_9_13;
  wire [`AWIDTH-1:0] c_addr_9_14;
  wire [`AWIDTH-1:0] c_addr_9_15;
  wire [`AWIDTH-1:0] c_addr_10_0;
  wire [`AWIDTH-1:0] c_addr_10_1;
  wire [`AWIDTH-1:0] c_addr_10_2;
  wire [`AWIDTH-1:0] c_addr_10_3;
  wire [`AWIDTH-1:0] c_addr_10_4;
  wire [`AWIDTH-1:0] c_addr_10_5;
  wire [`AWIDTH-1:0] c_addr_10_6;
  wire [`AWIDTH-1:0] c_addr_10_7;
  wire [`AWIDTH-1:0] c_addr_10_8;
  wire [`AWIDTH-1:0] c_addr_10_9;
  wire [`AWIDTH-1:0] c_addr_10_10;
  wire [`AWIDTH-1:0] c_addr_10_11;
  wire [`AWIDTH-1:0] c_addr_10_12;
  wire [`AWIDTH-1:0] c_addr_10_13;
  wire [`AWIDTH-1:0] c_addr_10_14;
  wire [`AWIDTH-1:0] c_addr_10_15;
  wire [`AWIDTH-1:0] c_addr_11_0;
  wire [`AWIDTH-1:0] c_addr_11_1;
  wire [`AWIDTH-1:0] c_addr_11_2;
  wire [`AWIDTH-1:0] c_addr_11_3;
  wire [`AWIDTH-1:0] c_addr_11_4;
  wire [`AWIDTH-1:0] c_addr_11_5;
  wire [`AWIDTH-1:0] c_addr_11_6;
  wire [`AWIDTH-1:0] c_addr_11_7;
  wire [`AWIDTH-1:0] c_addr_11_8;
  wire [`AWIDTH-1:0] c_addr_11_9;
  wire [`AWIDTH-1:0] c_addr_11_10;
  wire [`AWIDTH-1:0] c_addr_11_11;
  wire [`AWIDTH-1:0] c_addr_11_12;
  wire [`AWIDTH-1:0] c_addr_11_13;
  wire [`AWIDTH-1:0] c_addr_11_14;
  wire [`AWIDTH-1:0] c_addr_11_15;
  wire [`AWIDTH-1:0] c_addr_12_0;
  wire [`AWIDTH-1:0] c_addr_12_1;
  wire [`AWIDTH-1:0] c_addr_12_2;
  wire [`AWIDTH-1:0] c_addr_12_3;
  wire [`AWIDTH-1:0] c_addr_12_4;
  wire [`AWIDTH-1:0] c_addr_12_5;
  wire [`AWIDTH-1:0] c_addr_12_6;
  wire [`AWIDTH-1:0] c_addr_12_7;
  wire [`AWIDTH-1:0] c_addr_12_8;
  wire [`AWIDTH-1:0] c_addr_12_9;
  wire [`AWIDTH-1:0] c_addr_12_10;
  wire [`AWIDTH-1:0] c_addr_12_11;
  wire [`AWIDTH-1:0] c_addr_12_12;
  wire [`AWIDTH-1:0] c_addr_12_13;
  wire [`AWIDTH-1:0] c_addr_12_14;
  wire [`AWIDTH-1:0] c_addr_12_15;
  wire [`AWIDTH-1:0] c_addr_13_0;
  wire [`AWIDTH-1:0] c_addr_13_1;
  wire [`AWIDTH-1:0] c_addr_13_2;
  wire [`AWIDTH-1:0] c_addr_13_3;
  wire [`AWIDTH-1:0] c_addr_13_4;
  wire [`AWIDTH-1:0] c_addr_13_5;
  wire [`AWIDTH-1:0] c_addr_13_6;
  wire [`AWIDTH-1:0] c_addr_13_7;
  wire [`AWIDTH-1:0] c_addr_13_8;
  wire [`AWIDTH-1:0] c_addr_13_9;
  wire [`AWIDTH-1:0] c_addr_13_10;
  wire [`AWIDTH-1:0] c_addr_13_11;
  wire [`AWIDTH-1:0] c_addr_13_12;
  wire [`AWIDTH-1:0] c_addr_13_13;
  wire [`AWIDTH-1:0] c_addr_13_14;
  wire [`AWIDTH-1:0] c_addr_13_15;
  wire [`AWIDTH-1:0] c_addr_14_0;
  wire [`AWIDTH-1:0] c_addr_14_1;
  wire [`AWIDTH-1:0] c_addr_14_2;
  wire [`AWIDTH-1:0] c_addr_14_3;
  wire [`AWIDTH-1:0] c_addr_14_4;
  wire [`AWIDTH-1:0] c_addr_14_5;
  wire [`AWIDTH-1:0] c_addr_14_6;
  wire [`AWIDTH-1:0] c_addr_14_7;
  wire [`AWIDTH-1:0] c_addr_14_8;
  wire [`AWIDTH-1:0] c_addr_14_9;
  wire [`AWIDTH-1:0] c_addr_14_10;
  wire [`AWIDTH-1:0] c_addr_14_11;
  wire [`AWIDTH-1:0] c_addr_14_12;
  wire [`AWIDTH-1:0] c_addr_14_13;
  wire [`AWIDTH-1:0] c_addr_14_14;
  wire [`AWIDTH-1:0] c_addr_14_15;
  wire [`AWIDTH-1:0] c_addr_15_0;
  wire [`AWIDTH-1:0] c_addr_15_1;
  wire [`AWIDTH-1:0] c_addr_15_2;
  wire [`AWIDTH-1:0] c_addr_15_3;
  wire [`AWIDTH-1:0] c_addr_15_4;
  wire [`AWIDTH-1:0] c_addr_15_5;
  wire [`AWIDTH-1:0] c_addr_15_6;
  wire [`AWIDTH-1:0] c_addr_15_7;
  wire [`AWIDTH-1:0] c_addr_15_8;
  wire [`AWIDTH-1:0] c_addr_15_9;
  wire [`AWIDTH-1:0] c_addr_15_10;
  wire [`AWIDTH-1:0] c_addr_15_11;
  wire [`AWIDTH-1:0] c_addr_15_12;
  wire [`AWIDTH-1:0] c_addr_15_13;
  wire [`AWIDTH-1:0] c_addr_15_14;
  wire [`AWIDTH-1:0] c_addr_15_15;

  wire [`AWIDTH-1:0] c_addr_muxed_0_0;
  wire [`AWIDTH-1:0] c_addr_muxed_0_1;
  wire [`AWIDTH-1:0] c_addr_muxed_0_2;
  wire [`AWIDTH-1:0] c_addr_muxed_0_3;
  wire [`AWIDTH-1:0] c_addr_muxed_0_4;
  wire [`AWIDTH-1:0] c_addr_muxed_0_5;
  wire [`AWIDTH-1:0] c_addr_muxed_0_6;
  wire [`AWIDTH-1:0] c_addr_muxed_0_7;
  wire [`AWIDTH-1:0] c_addr_muxed_0_8;
  wire [`AWIDTH-1:0] c_addr_muxed_0_9;
  wire [`AWIDTH-1:0] c_addr_muxed_0_10;
  wire [`AWIDTH-1:0] c_addr_muxed_0_11;
  wire [`AWIDTH-1:0] c_addr_muxed_0_12;
  wire [`AWIDTH-1:0] c_addr_muxed_0_13;
  wire [`AWIDTH-1:0] c_addr_muxed_0_14;
  wire [`AWIDTH-1:0] c_addr_muxed_0_15;
  wire [`AWIDTH-1:0] c_addr_muxed_1_0;
  wire [`AWIDTH-1:0] c_addr_muxed_1_1;
  wire [`AWIDTH-1:0] c_addr_muxed_1_2;
  wire [`AWIDTH-1:0] c_addr_muxed_1_3;
  wire [`AWIDTH-1:0] c_addr_muxed_1_4;
  wire [`AWIDTH-1:0] c_addr_muxed_1_5;
  wire [`AWIDTH-1:0] c_addr_muxed_1_6;
  wire [`AWIDTH-1:0] c_addr_muxed_1_7;
  wire [`AWIDTH-1:0] c_addr_muxed_1_8;
  wire [`AWIDTH-1:0] c_addr_muxed_1_9;
  wire [`AWIDTH-1:0] c_addr_muxed_1_10;
  wire [`AWIDTH-1:0] c_addr_muxed_1_11;
  wire [`AWIDTH-1:0] c_addr_muxed_1_12;
  wire [`AWIDTH-1:0] c_addr_muxed_1_13;
  wire [`AWIDTH-1:0] c_addr_muxed_1_14;
  wire [`AWIDTH-1:0] c_addr_muxed_1_15;
  wire [`AWIDTH-1:0] c_addr_muxed_2_0;
  wire [`AWIDTH-1:0] c_addr_muxed_2_1;
  wire [`AWIDTH-1:0] c_addr_muxed_2_2;
  wire [`AWIDTH-1:0] c_addr_muxed_2_3;
  wire [`AWIDTH-1:0] c_addr_muxed_2_4;
  wire [`AWIDTH-1:0] c_addr_muxed_2_5;
  wire [`AWIDTH-1:0] c_addr_muxed_2_6;
  wire [`AWIDTH-1:0] c_addr_muxed_2_7;
  wire [`AWIDTH-1:0] c_addr_muxed_2_8;
  wire [`AWIDTH-1:0] c_addr_muxed_2_9;
  wire [`AWIDTH-1:0] c_addr_muxed_2_10;
  wire [`AWIDTH-1:0] c_addr_muxed_2_11;
  wire [`AWIDTH-1:0] c_addr_muxed_2_12;
  wire [`AWIDTH-1:0] c_addr_muxed_2_13;
  wire [`AWIDTH-1:0] c_addr_muxed_2_14;
  wire [`AWIDTH-1:0] c_addr_muxed_2_15;
  wire [`AWIDTH-1:0] c_addr_muxed_3_0;
  wire [`AWIDTH-1:0] c_addr_muxed_3_1;
  wire [`AWIDTH-1:0] c_addr_muxed_3_2;
  wire [`AWIDTH-1:0] c_addr_muxed_3_3;
  wire [`AWIDTH-1:0] c_addr_muxed_3_4;
  wire [`AWIDTH-1:0] c_addr_muxed_3_5;
  wire [`AWIDTH-1:0] c_addr_muxed_3_6;
  wire [`AWIDTH-1:0] c_addr_muxed_3_7;
  wire [`AWIDTH-1:0] c_addr_muxed_3_8;
  wire [`AWIDTH-1:0] c_addr_muxed_3_9;
  wire [`AWIDTH-1:0] c_addr_muxed_3_10;
  wire [`AWIDTH-1:0] c_addr_muxed_3_11;
  wire [`AWIDTH-1:0] c_addr_muxed_3_12;
  wire [`AWIDTH-1:0] c_addr_muxed_3_13;
  wire [`AWIDTH-1:0] c_addr_muxed_3_14;
  wire [`AWIDTH-1:0] c_addr_muxed_3_15;
  wire [`AWIDTH-1:0] c_addr_muxed_4_0;
  wire [`AWIDTH-1:0] c_addr_muxed_4_1;
  wire [`AWIDTH-1:0] c_addr_muxed_4_2;
  wire [`AWIDTH-1:0] c_addr_muxed_4_3;
  wire [`AWIDTH-1:0] c_addr_muxed_4_4;
  wire [`AWIDTH-1:0] c_addr_muxed_4_5;
  wire [`AWIDTH-1:0] c_addr_muxed_4_6;
  wire [`AWIDTH-1:0] c_addr_muxed_4_7;
  wire [`AWIDTH-1:0] c_addr_muxed_4_8;
  wire [`AWIDTH-1:0] c_addr_muxed_4_9;
  wire [`AWIDTH-1:0] c_addr_muxed_4_10;
  wire [`AWIDTH-1:0] c_addr_muxed_4_11;
  wire [`AWIDTH-1:0] c_addr_muxed_4_12;
  wire [`AWIDTH-1:0] c_addr_muxed_4_13;
  wire [`AWIDTH-1:0] c_addr_muxed_4_14;
  wire [`AWIDTH-1:0] c_addr_muxed_4_15;
  wire [`AWIDTH-1:0] c_addr_muxed_5_0;
  wire [`AWIDTH-1:0] c_addr_muxed_5_1;
  wire [`AWIDTH-1:0] c_addr_muxed_5_2;
  wire [`AWIDTH-1:0] c_addr_muxed_5_3;
  wire [`AWIDTH-1:0] c_addr_muxed_5_4;
  wire [`AWIDTH-1:0] c_addr_muxed_5_5;
  wire [`AWIDTH-1:0] c_addr_muxed_5_6;
  wire [`AWIDTH-1:0] c_addr_muxed_5_7;
  wire [`AWIDTH-1:0] c_addr_muxed_5_8;
  wire [`AWIDTH-1:0] c_addr_muxed_5_9;
  wire [`AWIDTH-1:0] c_addr_muxed_5_10;
  wire [`AWIDTH-1:0] c_addr_muxed_5_11;
  wire [`AWIDTH-1:0] c_addr_muxed_5_12;
  wire [`AWIDTH-1:0] c_addr_muxed_5_13;
  wire [`AWIDTH-1:0] c_addr_muxed_5_14;
  wire [`AWIDTH-1:0] c_addr_muxed_5_15;
  wire [`AWIDTH-1:0] c_addr_muxed_6_0;
  wire [`AWIDTH-1:0] c_addr_muxed_6_1;
  wire [`AWIDTH-1:0] c_addr_muxed_6_2;
  wire [`AWIDTH-1:0] c_addr_muxed_6_3;
  wire [`AWIDTH-1:0] c_addr_muxed_6_4;
  wire [`AWIDTH-1:0] c_addr_muxed_6_5;
  wire [`AWIDTH-1:0] c_addr_muxed_6_6;
  wire [`AWIDTH-1:0] c_addr_muxed_6_7;
  wire [`AWIDTH-1:0] c_addr_muxed_6_8;
  wire [`AWIDTH-1:0] c_addr_muxed_6_9;
  wire [`AWIDTH-1:0] c_addr_muxed_6_10;
  wire [`AWIDTH-1:0] c_addr_muxed_6_11;
  wire [`AWIDTH-1:0] c_addr_muxed_6_12;
  wire [`AWIDTH-1:0] c_addr_muxed_6_13;
  wire [`AWIDTH-1:0] c_addr_muxed_6_14;
  wire [`AWIDTH-1:0] c_addr_muxed_6_15;
  wire [`AWIDTH-1:0] c_addr_muxed_7_0;
  wire [`AWIDTH-1:0] c_addr_muxed_7_1;
  wire [`AWIDTH-1:0] c_addr_muxed_7_2;
  wire [`AWIDTH-1:0] c_addr_muxed_7_3;
  wire [`AWIDTH-1:0] c_addr_muxed_7_4;
  wire [`AWIDTH-1:0] c_addr_muxed_7_5;
  wire [`AWIDTH-1:0] c_addr_muxed_7_6;
  wire [`AWIDTH-1:0] c_addr_muxed_7_7;
  wire [`AWIDTH-1:0] c_addr_muxed_7_8;
  wire [`AWIDTH-1:0] c_addr_muxed_7_9;
  wire [`AWIDTH-1:0] c_addr_muxed_7_10;
  wire [`AWIDTH-1:0] c_addr_muxed_7_11;
  wire [`AWIDTH-1:0] c_addr_muxed_7_12;
  wire [`AWIDTH-1:0] c_addr_muxed_7_13;
  wire [`AWIDTH-1:0] c_addr_muxed_7_14;
  wire [`AWIDTH-1:0] c_addr_muxed_7_15;
  wire [`AWIDTH-1:0] c_addr_muxed_8_0;
  wire [`AWIDTH-1:0] c_addr_muxed_8_1;
  wire [`AWIDTH-1:0] c_addr_muxed_8_2;
  wire [`AWIDTH-1:0] c_addr_muxed_8_3;
  wire [`AWIDTH-1:0] c_addr_muxed_8_4;
  wire [`AWIDTH-1:0] c_addr_muxed_8_5;
  wire [`AWIDTH-1:0] c_addr_muxed_8_6;
  wire [`AWIDTH-1:0] c_addr_muxed_8_7;
  wire [`AWIDTH-1:0] c_addr_muxed_8_8;
  wire [`AWIDTH-1:0] c_addr_muxed_8_9;
  wire [`AWIDTH-1:0] c_addr_muxed_8_10;
  wire [`AWIDTH-1:0] c_addr_muxed_8_11;
  wire [`AWIDTH-1:0] c_addr_muxed_8_12;
  wire [`AWIDTH-1:0] c_addr_muxed_8_13;
  wire [`AWIDTH-1:0] c_addr_muxed_8_14;
  wire [`AWIDTH-1:0] c_addr_muxed_8_15;
  wire [`AWIDTH-1:0] c_addr_muxed_9_0;
  wire [`AWIDTH-1:0] c_addr_muxed_9_1;
  wire [`AWIDTH-1:0] c_addr_muxed_9_2;
  wire [`AWIDTH-1:0] c_addr_muxed_9_3;
  wire [`AWIDTH-1:0] c_addr_muxed_9_4;
  wire [`AWIDTH-1:0] c_addr_muxed_9_5;
  wire [`AWIDTH-1:0] c_addr_muxed_9_6;
  wire [`AWIDTH-1:0] c_addr_muxed_9_7;
  wire [`AWIDTH-1:0] c_addr_muxed_9_8;
  wire [`AWIDTH-1:0] c_addr_muxed_9_9;
  wire [`AWIDTH-1:0] c_addr_muxed_9_10;
  wire [`AWIDTH-1:0] c_addr_muxed_9_11;
  wire [`AWIDTH-1:0] c_addr_muxed_9_12;
  wire [`AWIDTH-1:0] c_addr_muxed_9_13;
  wire [`AWIDTH-1:0] c_addr_muxed_9_14;
  wire [`AWIDTH-1:0] c_addr_muxed_9_15;
  wire [`AWIDTH-1:0] c_addr_muxed_10_0;
  wire [`AWIDTH-1:0] c_addr_muxed_10_1;
  wire [`AWIDTH-1:0] c_addr_muxed_10_2;
  wire [`AWIDTH-1:0] c_addr_muxed_10_3;
  wire [`AWIDTH-1:0] c_addr_muxed_10_4;
  wire [`AWIDTH-1:0] c_addr_muxed_10_5;
  wire [`AWIDTH-1:0] c_addr_muxed_10_6;
  wire [`AWIDTH-1:0] c_addr_muxed_10_7;
  wire [`AWIDTH-1:0] c_addr_muxed_10_8;
  wire [`AWIDTH-1:0] c_addr_muxed_10_9;
  wire [`AWIDTH-1:0] c_addr_muxed_10_10;
  wire [`AWIDTH-1:0] c_addr_muxed_10_11;
  wire [`AWIDTH-1:0] c_addr_muxed_10_12;
  wire [`AWIDTH-1:0] c_addr_muxed_10_13;
  wire [`AWIDTH-1:0] c_addr_muxed_10_14;
  wire [`AWIDTH-1:0] c_addr_muxed_10_15;
  wire [`AWIDTH-1:0] c_addr_muxed_11_0;
  wire [`AWIDTH-1:0] c_addr_muxed_11_1;
  wire [`AWIDTH-1:0] c_addr_muxed_11_2;
  wire [`AWIDTH-1:0] c_addr_muxed_11_3;
  wire [`AWIDTH-1:0] c_addr_muxed_11_4;
  wire [`AWIDTH-1:0] c_addr_muxed_11_5;
  wire [`AWIDTH-1:0] c_addr_muxed_11_6;
  wire [`AWIDTH-1:0] c_addr_muxed_11_7;
  wire [`AWIDTH-1:0] c_addr_muxed_11_8;
  wire [`AWIDTH-1:0] c_addr_muxed_11_9;
  wire [`AWIDTH-1:0] c_addr_muxed_11_10;
  wire [`AWIDTH-1:0] c_addr_muxed_11_11;
  wire [`AWIDTH-1:0] c_addr_muxed_11_12;
  wire [`AWIDTH-1:0] c_addr_muxed_11_13;
  wire [`AWIDTH-1:0] c_addr_muxed_11_14;
  wire [`AWIDTH-1:0] c_addr_muxed_11_15;
  wire [`AWIDTH-1:0] c_addr_muxed_12_0;
  wire [`AWIDTH-1:0] c_addr_muxed_12_1;
  wire [`AWIDTH-1:0] c_addr_muxed_12_2;
  wire [`AWIDTH-1:0] c_addr_muxed_12_3;
  wire [`AWIDTH-1:0] c_addr_muxed_12_4;
  wire [`AWIDTH-1:0] c_addr_muxed_12_5;
  wire [`AWIDTH-1:0] c_addr_muxed_12_6;
  wire [`AWIDTH-1:0] c_addr_muxed_12_7;
  wire [`AWIDTH-1:0] c_addr_muxed_12_8;
  wire [`AWIDTH-1:0] c_addr_muxed_12_9;
  wire [`AWIDTH-1:0] c_addr_muxed_12_10;
  wire [`AWIDTH-1:0] c_addr_muxed_12_11;
  wire [`AWIDTH-1:0] c_addr_muxed_12_12;
  wire [`AWIDTH-1:0] c_addr_muxed_12_13;
  wire [`AWIDTH-1:0] c_addr_muxed_12_14;
  wire [`AWIDTH-1:0] c_addr_muxed_12_15;
  wire [`AWIDTH-1:0] c_addr_muxed_13_0;
  wire [`AWIDTH-1:0] c_addr_muxed_13_1;
  wire [`AWIDTH-1:0] c_addr_muxed_13_2;
  wire [`AWIDTH-1:0] c_addr_muxed_13_3;
  wire [`AWIDTH-1:0] c_addr_muxed_13_4;
  wire [`AWIDTH-1:0] c_addr_muxed_13_5;
  wire [`AWIDTH-1:0] c_addr_muxed_13_6;
  wire [`AWIDTH-1:0] c_addr_muxed_13_7;
  wire [`AWIDTH-1:0] c_addr_muxed_13_8;
  wire [`AWIDTH-1:0] c_addr_muxed_13_9;
  wire [`AWIDTH-1:0] c_addr_muxed_13_10;
  wire [`AWIDTH-1:0] c_addr_muxed_13_11;
  wire [`AWIDTH-1:0] c_addr_muxed_13_12;
  wire [`AWIDTH-1:0] c_addr_muxed_13_13;
  wire [`AWIDTH-1:0] c_addr_muxed_13_14;
  wire [`AWIDTH-1:0] c_addr_muxed_13_15;
  wire [`AWIDTH-1:0] c_addr_muxed_14_0;
  wire [`AWIDTH-1:0] c_addr_muxed_14_1;
  wire [`AWIDTH-1:0] c_addr_muxed_14_2;
  wire [`AWIDTH-1:0] c_addr_muxed_14_3;
  wire [`AWIDTH-1:0] c_addr_muxed_14_4;
  wire [`AWIDTH-1:0] c_addr_muxed_14_5;
  wire [`AWIDTH-1:0] c_addr_muxed_14_6;
  wire [`AWIDTH-1:0] c_addr_muxed_14_7;
  wire [`AWIDTH-1:0] c_addr_muxed_14_8;
  wire [`AWIDTH-1:0] c_addr_muxed_14_9;
  wire [`AWIDTH-1:0] c_addr_muxed_14_10;
  wire [`AWIDTH-1:0] c_addr_muxed_14_11;
  wire [`AWIDTH-1:0] c_addr_muxed_14_12;
  wire [`AWIDTH-1:0] c_addr_muxed_14_13;
  wire [`AWIDTH-1:0] c_addr_muxed_14_14;
  wire [`AWIDTH-1:0] c_addr_muxed_14_15;
  wire [`AWIDTH-1:0] c_addr_muxed_15_0;
  wire [`AWIDTH-1:0] c_addr_muxed_15_1;
  wire [`AWIDTH-1:0] c_addr_muxed_15_2;
  wire [`AWIDTH-1:0] c_addr_muxed_15_3;
  wire [`AWIDTH-1:0] c_addr_muxed_15_4;
  wire [`AWIDTH-1:0] c_addr_muxed_15_5;
  wire [`AWIDTH-1:0] c_addr_muxed_15_6;
  wire [`AWIDTH-1:0] c_addr_muxed_15_7;
  wire [`AWIDTH-1:0] c_addr_muxed_15_8;
  wire [`AWIDTH-1:0] c_addr_muxed_15_9;
  wire [`AWIDTH-1:0] c_addr_muxed_15_10;
  wire [`AWIDTH-1:0] c_addr_muxed_15_11;
  wire [`AWIDTH-1:0] c_addr_muxed_15_12;
  wire [`AWIDTH-1:0] c_addr_muxed_15_13;
  wire [`AWIDTH-1:0] c_addr_muxed_15_14;
  wire [`AWIDTH-1:0] c_addr_muxed_15_15;

  reg [`AWIDTH-1:0] c_addr_0_0_reg;
  reg [`AWIDTH-1:0] c_addr_0_1_reg;
  reg [`AWIDTH-1:0] c_addr_0_2_reg;
  reg [`AWIDTH-1:0] c_addr_0_3_reg;
  reg [`AWIDTH-1:0] c_addr_0_4_reg;
  reg [`AWIDTH-1:0] c_addr_0_5_reg;
  reg [`AWIDTH-1:0] c_addr_0_6_reg;
  reg [`AWIDTH-1:0] c_addr_0_7_reg;
  reg [`AWIDTH-1:0] c_addr_0_8_reg;
  reg [`AWIDTH-1:0] c_addr_0_9_reg;
  reg [`AWIDTH-1:0] c_addr_0_10_reg;
  reg [`AWIDTH-1:0] c_addr_0_11_reg;
  reg [`AWIDTH-1:0] c_addr_0_12_reg;
  reg [`AWIDTH-1:0] c_addr_0_13_reg;
  reg [`AWIDTH-1:0] c_addr_0_14_reg;
  reg [`AWIDTH-1:0] c_addr_0_15_reg;
  reg [`AWIDTH-1:0] c_addr_1_0_reg;
  reg [`AWIDTH-1:0] c_addr_1_1_reg;
  reg [`AWIDTH-1:0] c_addr_1_2_reg;
  reg [`AWIDTH-1:0] c_addr_1_3_reg;
  reg [`AWIDTH-1:0] c_addr_1_4_reg;
  reg [`AWIDTH-1:0] c_addr_1_5_reg;
  reg [`AWIDTH-1:0] c_addr_1_6_reg;
  reg [`AWIDTH-1:0] c_addr_1_7_reg;
  reg [`AWIDTH-1:0] c_addr_1_8_reg;
  reg [`AWIDTH-1:0] c_addr_1_9_reg;
  reg [`AWIDTH-1:0] c_addr_1_10_reg;
  reg [`AWIDTH-1:0] c_addr_1_11_reg;
  reg [`AWIDTH-1:0] c_addr_1_12_reg;
  reg [`AWIDTH-1:0] c_addr_1_13_reg;
  reg [`AWIDTH-1:0] c_addr_1_14_reg;
  reg [`AWIDTH-1:0] c_addr_1_15_reg;
  reg [`AWIDTH-1:0] c_addr_2_0_reg;
  reg [`AWIDTH-1:0] c_addr_2_1_reg;
  reg [`AWIDTH-1:0] c_addr_2_2_reg;
  reg [`AWIDTH-1:0] c_addr_2_3_reg;
  reg [`AWIDTH-1:0] c_addr_2_4_reg;
  reg [`AWIDTH-1:0] c_addr_2_5_reg;
  reg [`AWIDTH-1:0] c_addr_2_6_reg;
  reg [`AWIDTH-1:0] c_addr_2_7_reg;
  reg [`AWIDTH-1:0] c_addr_2_8_reg;
  reg [`AWIDTH-1:0] c_addr_2_9_reg;
  reg [`AWIDTH-1:0] c_addr_2_10_reg;
  reg [`AWIDTH-1:0] c_addr_2_11_reg;
  reg [`AWIDTH-1:0] c_addr_2_12_reg;
  reg [`AWIDTH-1:0] c_addr_2_13_reg;
  reg [`AWIDTH-1:0] c_addr_2_14_reg;
  reg [`AWIDTH-1:0] c_addr_2_15_reg;
  reg [`AWIDTH-1:0] c_addr_3_0_reg;
  reg [`AWIDTH-1:0] c_addr_3_1_reg;
  reg [`AWIDTH-1:0] c_addr_3_2_reg;
  reg [`AWIDTH-1:0] c_addr_3_3_reg;
  reg [`AWIDTH-1:0] c_addr_3_4_reg;
  reg [`AWIDTH-1:0] c_addr_3_5_reg;
  reg [`AWIDTH-1:0] c_addr_3_6_reg;
  reg [`AWIDTH-1:0] c_addr_3_7_reg;
  reg [`AWIDTH-1:0] c_addr_3_8_reg;
  reg [`AWIDTH-1:0] c_addr_3_9_reg;
  reg [`AWIDTH-1:0] c_addr_3_10_reg;
  reg [`AWIDTH-1:0] c_addr_3_11_reg;
  reg [`AWIDTH-1:0] c_addr_3_12_reg;
  reg [`AWIDTH-1:0] c_addr_3_13_reg;
  reg [`AWIDTH-1:0] c_addr_3_14_reg;
  reg [`AWIDTH-1:0] c_addr_3_15_reg;
  reg [`AWIDTH-1:0] c_addr_4_0_reg;
  reg [`AWIDTH-1:0] c_addr_4_1_reg;
  reg [`AWIDTH-1:0] c_addr_4_2_reg;
  reg [`AWIDTH-1:0] c_addr_4_3_reg;
  reg [`AWIDTH-1:0] c_addr_4_4_reg;
  reg [`AWIDTH-1:0] c_addr_4_5_reg;
  reg [`AWIDTH-1:0] c_addr_4_6_reg;
  reg [`AWIDTH-1:0] c_addr_4_7_reg;
  reg [`AWIDTH-1:0] c_addr_4_8_reg;
  reg [`AWIDTH-1:0] c_addr_4_9_reg;
  reg [`AWIDTH-1:0] c_addr_4_10_reg;
  reg [`AWIDTH-1:0] c_addr_4_11_reg;
  reg [`AWIDTH-1:0] c_addr_4_12_reg;
  reg [`AWIDTH-1:0] c_addr_4_13_reg;
  reg [`AWIDTH-1:0] c_addr_4_14_reg;
  reg [`AWIDTH-1:0] c_addr_4_15_reg;
  reg [`AWIDTH-1:0] c_addr_5_0_reg;
  reg [`AWIDTH-1:0] c_addr_5_1_reg;
  reg [`AWIDTH-1:0] c_addr_5_2_reg;
  reg [`AWIDTH-1:0] c_addr_5_3_reg;
  reg [`AWIDTH-1:0] c_addr_5_4_reg;
  reg [`AWIDTH-1:0] c_addr_5_5_reg;
  reg [`AWIDTH-1:0] c_addr_5_6_reg;
  reg [`AWIDTH-1:0] c_addr_5_7_reg;
  reg [`AWIDTH-1:0] c_addr_5_8_reg;
  reg [`AWIDTH-1:0] c_addr_5_9_reg;
  reg [`AWIDTH-1:0] c_addr_5_10_reg;
  reg [`AWIDTH-1:0] c_addr_5_11_reg;
  reg [`AWIDTH-1:0] c_addr_5_12_reg;
  reg [`AWIDTH-1:0] c_addr_5_13_reg;
  reg [`AWIDTH-1:0] c_addr_5_14_reg;
  reg [`AWIDTH-1:0] c_addr_5_15_reg;
  reg [`AWIDTH-1:0] c_addr_6_0_reg;
  reg [`AWIDTH-1:0] c_addr_6_1_reg;
  reg [`AWIDTH-1:0] c_addr_6_2_reg;
  reg [`AWIDTH-1:0] c_addr_6_3_reg;
  reg [`AWIDTH-1:0] c_addr_6_4_reg;
  reg [`AWIDTH-1:0] c_addr_6_5_reg;
  reg [`AWIDTH-1:0] c_addr_6_6_reg;
  reg [`AWIDTH-1:0] c_addr_6_7_reg;
  reg [`AWIDTH-1:0] c_addr_6_8_reg;
  reg [`AWIDTH-1:0] c_addr_6_9_reg;
  reg [`AWIDTH-1:0] c_addr_6_10_reg;
  reg [`AWIDTH-1:0] c_addr_6_11_reg;
  reg [`AWIDTH-1:0] c_addr_6_12_reg;
  reg [`AWIDTH-1:0] c_addr_6_13_reg;
  reg [`AWIDTH-1:0] c_addr_6_14_reg;
  reg [`AWIDTH-1:0] c_addr_6_15_reg;
  reg [`AWIDTH-1:0] c_addr_7_0_reg;
  reg [`AWIDTH-1:0] c_addr_7_1_reg;
  reg [`AWIDTH-1:0] c_addr_7_2_reg;
  reg [`AWIDTH-1:0] c_addr_7_3_reg;
  reg [`AWIDTH-1:0] c_addr_7_4_reg;
  reg [`AWIDTH-1:0] c_addr_7_5_reg;
  reg [`AWIDTH-1:0] c_addr_7_6_reg;
  reg [`AWIDTH-1:0] c_addr_7_7_reg;
  reg [`AWIDTH-1:0] c_addr_7_8_reg;
  reg [`AWIDTH-1:0] c_addr_7_9_reg;
  reg [`AWIDTH-1:0] c_addr_7_10_reg;
  reg [`AWIDTH-1:0] c_addr_7_11_reg;
  reg [`AWIDTH-1:0] c_addr_7_12_reg;
  reg [`AWIDTH-1:0] c_addr_7_13_reg;
  reg [`AWIDTH-1:0] c_addr_7_14_reg;
  reg [`AWIDTH-1:0] c_addr_7_15_reg;
  reg [`AWIDTH-1:0] c_addr_8_0_reg;
  reg [`AWIDTH-1:0] c_addr_8_1_reg;
  reg [`AWIDTH-1:0] c_addr_8_2_reg;
  reg [`AWIDTH-1:0] c_addr_8_3_reg;
  reg [`AWIDTH-1:0] c_addr_8_4_reg;
  reg [`AWIDTH-1:0] c_addr_8_5_reg;
  reg [`AWIDTH-1:0] c_addr_8_6_reg;
  reg [`AWIDTH-1:0] c_addr_8_7_reg;
  reg [`AWIDTH-1:0] c_addr_8_8_reg;
  reg [`AWIDTH-1:0] c_addr_8_9_reg;
  reg [`AWIDTH-1:0] c_addr_8_10_reg;
  reg [`AWIDTH-1:0] c_addr_8_11_reg;
  reg [`AWIDTH-1:0] c_addr_8_12_reg;
  reg [`AWIDTH-1:0] c_addr_8_13_reg;
  reg [`AWIDTH-1:0] c_addr_8_14_reg;
  reg [`AWIDTH-1:0] c_addr_8_15_reg;
  reg [`AWIDTH-1:0] c_addr_9_0_reg;
  reg [`AWIDTH-1:0] c_addr_9_1_reg;
  reg [`AWIDTH-1:0] c_addr_9_2_reg;
  reg [`AWIDTH-1:0] c_addr_9_3_reg;
  reg [`AWIDTH-1:0] c_addr_9_4_reg;
  reg [`AWIDTH-1:0] c_addr_9_5_reg;
  reg [`AWIDTH-1:0] c_addr_9_6_reg;
  reg [`AWIDTH-1:0] c_addr_9_7_reg;
  reg [`AWIDTH-1:0] c_addr_9_8_reg;
  reg [`AWIDTH-1:0] c_addr_9_9_reg;
  reg [`AWIDTH-1:0] c_addr_9_10_reg;
  reg [`AWIDTH-1:0] c_addr_9_11_reg;
  reg [`AWIDTH-1:0] c_addr_9_12_reg;
  reg [`AWIDTH-1:0] c_addr_9_13_reg;
  reg [`AWIDTH-1:0] c_addr_9_14_reg;
  reg [`AWIDTH-1:0] c_addr_9_15_reg;
  reg [`AWIDTH-1:0] c_addr_10_0_reg;
  reg [`AWIDTH-1:0] c_addr_10_1_reg;
  reg [`AWIDTH-1:0] c_addr_10_2_reg;
  reg [`AWIDTH-1:0] c_addr_10_3_reg;
  reg [`AWIDTH-1:0] c_addr_10_4_reg;
  reg [`AWIDTH-1:0] c_addr_10_5_reg;
  reg [`AWIDTH-1:0] c_addr_10_6_reg;
  reg [`AWIDTH-1:0] c_addr_10_7_reg;
  reg [`AWIDTH-1:0] c_addr_10_8_reg;
  reg [`AWIDTH-1:0] c_addr_10_9_reg;
  reg [`AWIDTH-1:0] c_addr_10_10_reg;
  reg [`AWIDTH-1:0] c_addr_10_11_reg;
  reg [`AWIDTH-1:0] c_addr_10_12_reg;
  reg [`AWIDTH-1:0] c_addr_10_13_reg;
  reg [`AWIDTH-1:0] c_addr_10_14_reg;
  reg [`AWIDTH-1:0] c_addr_10_15_reg;
  reg [`AWIDTH-1:0] c_addr_11_0_reg;
  reg [`AWIDTH-1:0] c_addr_11_1_reg;
  reg [`AWIDTH-1:0] c_addr_11_2_reg;
  reg [`AWIDTH-1:0] c_addr_11_3_reg;
  reg [`AWIDTH-1:0] c_addr_11_4_reg;
  reg [`AWIDTH-1:0] c_addr_11_5_reg;
  reg [`AWIDTH-1:0] c_addr_11_6_reg;
  reg [`AWIDTH-1:0] c_addr_11_7_reg;
  reg [`AWIDTH-1:0] c_addr_11_8_reg;
  reg [`AWIDTH-1:0] c_addr_11_9_reg;
  reg [`AWIDTH-1:0] c_addr_11_10_reg;
  reg [`AWIDTH-1:0] c_addr_11_11_reg;
  reg [`AWIDTH-1:0] c_addr_11_12_reg;
  reg [`AWIDTH-1:0] c_addr_11_13_reg;
  reg [`AWIDTH-1:0] c_addr_11_14_reg;
  reg [`AWIDTH-1:0] c_addr_11_15_reg;
  reg [`AWIDTH-1:0] c_addr_12_0_reg;
  reg [`AWIDTH-1:0] c_addr_12_1_reg;
  reg [`AWIDTH-1:0] c_addr_12_2_reg;
  reg [`AWIDTH-1:0] c_addr_12_3_reg;
  reg [`AWIDTH-1:0] c_addr_12_4_reg;
  reg [`AWIDTH-1:0] c_addr_12_5_reg;
  reg [`AWIDTH-1:0] c_addr_12_6_reg;
  reg [`AWIDTH-1:0] c_addr_12_7_reg;
  reg [`AWIDTH-1:0] c_addr_12_8_reg;
  reg [`AWIDTH-1:0] c_addr_12_9_reg;
  reg [`AWIDTH-1:0] c_addr_12_10_reg;
  reg [`AWIDTH-1:0] c_addr_12_11_reg;
  reg [`AWIDTH-1:0] c_addr_12_12_reg;
  reg [`AWIDTH-1:0] c_addr_12_13_reg;
  reg [`AWIDTH-1:0] c_addr_12_14_reg;
  reg [`AWIDTH-1:0] c_addr_12_15_reg;
  reg [`AWIDTH-1:0] c_addr_13_0_reg;
  reg [`AWIDTH-1:0] c_addr_13_1_reg;
  reg [`AWIDTH-1:0] c_addr_13_2_reg;
  reg [`AWIDTH-1:0] c_addr_13_3_reg;
  reg [`AWIDTH-1:0] c_addr_13_4_reg;
  reg [`AWIDTH-1:0] c_addr_13_5_reg;
  reg [`AWIDTH-1:0] c_addr_13_6_reg;
  reg [`AWIDTH-1:0] c_addr_13_7_reg;
  reg [`AWIDTH-1:0] c_addr_13_8_reg;
  reg [`AWIDTH-1:0] c_addr_13_9_reg;
  reg [`AWIDTH-1:0] c_addr_13_10_reg;
  reg [`AWIDTH-1:0] c_addr_13_11_reg;
  reg [`AWIDTH-1:0] c_addr_13_12_reg;
  reg [`AWIDTH-1:0] c_addr_13_13_reg;
  reg [`AWIDTH-1:0] c_addr_13_14_reg;
  reg [`AWIDTH-1:0] c_addr_13_15_reg;
  reg [`AWIDTH-1:0] c_addr_14_0_reg;
  reg [`AWIDTH-1:0] c_addr_14_1_reg;
  reg [`AWIDTH-1:0] c_addr_14_2_reg;
  reg [`AWIDTH-1:0] c_addr_14_3_reg;
  reg [`AWIDTH-1:0] c_addr_14_4_reg;
  reg [`AWIDTH-1:0] c_addr_14_5_reg;
  reg [`AWIDTH-1:0] c_addr_14_6_reg;
  reg [`AWIDTH-1:0] c_addr_14_7_reg;
  reg [`AWIDTH-1:0] c_addr_14_8_reg;
  reg [`AWIDTH-1:0] c_addr_14_9_reg;
  reg [`AWIDTH-1:0] c_addr_14_10_reg;
  reg [`AWIDTH-1:0] c_addr_14_11_reg;
  reg [`AWIDTH-1:0] c_addr_14_12_reg;
  reg [`AWIDTH-1:0] c_addr_14_13_reg;
  reg [`AWIDTH-1:0] c_addr_14_14_reg;
  reg [`AWIDTH-1:0] c_addr_14_15_reg;
  reg [`AWIDTH-1:0] c_addr_15_0_reg;
  reg [`AWIDTH-1:0] c_addr_15_1_reg;
  reg [`AWIDTH-1:0] c_addr_15_2_reg;
  reg [`AWIDTH-1:0] c_addr_15_3_reg;
  reg [`AWIDTH-1:0] c_addr_15_4_reg;
  reg [`AWIDTH-1:0] c_addr_15_5_reg;
  reg [`AWIDTH-1:0] c_addr_15_6_reg;
  reg [`AWIDTH-1:0] c_addr_15_7_reg;
  reg [`AWIDTH-1:0] c_addr_15_8_reg;
  reg [`AWIDTH-1:0] c_addr_15_9_reg;
  reg [`AWIDTH-1:0] c_addr_15_10_reg;
  reg [`AWIDTH-1:0] c_addr_15_11_reg;
  reg [`AWIDTH-1:0] c_addr_15_12_reg;
  reg [`AWIDTH-1:0] c_addr_15_13_reg;
  reg [`AWIDTH-1:0] c_addr_15_14_reg;
  reg [`AWIDTH-1:0] c_addr_15_15_reg;

  reg [`AWIDTH-1:0] c_addr_muxed_0_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_0_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_1_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_2_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_3_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_4_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_5_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_6_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_7_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_8_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_9_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_10_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_11_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_12_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_13_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_14_15_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_0_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_1_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_2_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_3_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_4_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_5_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_6_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_7_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_8_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_9_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_10_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_11_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_12_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_13_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_14_reg;
  reg [`AWIDTH-1:0] c_addr_muxed_15_15_reg;

  assign c_addr_muxed_0_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_0_reg;
  assign c_addr_muxed_0_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_1_reg;
  assign c_addr_muxed_0_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_2_reg;
  assign c_addr_muxed_0_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_3_reg;
  assign c_addr_muxed_0_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_4_reg;
  assign c_addr_muxed_0_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_5_reg;
  assign c_addr_muxed_0_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_6_reg;
  assign c_addr_muxed_0_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_7_reg;
  assign c_addr_muxed_0_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_8_reg;
  assign c_addr_muxed_0_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_9_reg;
  assign c_addr_muxed_0_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_10_reg;
  assign c_addr_muxed_0_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_11_reg;
  assign c_addr_muxed_0_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_12_reg;
  assign c_addr_muxed_0_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_13_reg;
  assign c_addr_muxed_0_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_14_reg;
  assign c_addr_muxed_0_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_0_15_reg;
  assign c_addr_muxed_1_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_0_reg;
  assign c_addr_muxed_1_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_1_reg;
  assign c_addr_muxed_1_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_2_reg;
  assign c_addr_muxed_1_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_3_reg;
  assign c_addr_muxed_1_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_4_reg;
  assign c_addr_muxed_1_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_5_reg;
  assign c_addr_muxed_1_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_6_reg;
  assign c_addr_muxed_1_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_7_reg;
  assign c_addr_muxed_1_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_8_reg;
  assign c_addr_muxed_1_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_9_reg;
  assign c_addr_muxed_1_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_10_reg;
  assign c_addr_muxed_1_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_11_reg;
  assign c_addr_muxed_1_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_12_reg;
  assign c_addr_muxed_1_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_13_reg;
  assign c_addr_muxed_1_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_14_reg;
  assign c_addr_muxed_1_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_1_15_reg;
  assign c_addr_muxed_2_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_0_reg;
  assign c_addr_muxed_2_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_1_reg;
  assign c_addr_muxed_2_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_2_reg;
  assign c_addr_muxed_2_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_3_reg;
  assign c_addr_muxed_2_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_4_reg;
  assign c_addr_muxed_2_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_5_reg;
  assign c_addr_muxed_2_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_6_reg;
  assign c_addr_muxed_2_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_7_reg;
  assign c_addr_muxed_2_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_8_reg;
  assign c_addr_muxed_2_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_9_reg;
  assign c_addr_muxed_2_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_10_reg;
  assign c_addr_muxed_2_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_11_reg;
  assign c_addr_muxed_2_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_12_reg;
  assign c_addr_muxed_2_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_13_reg;
  assign c_addr_muxed_2_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_14_reg;
  assign c_addr_muxed_2_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_2_15_reg;
  assign c_addr_muxed_3_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_0_reg;
  assign c_addr_muxed_3_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_1_reg;
  assign c_addr_muxed_3_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_2_reg;
  assign c_addr_muxed_3_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_3_reg;
  assign c_addr_muxed_3_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_4_reg;
  assign c_addr_muxed_3_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_5_reg;
  assign c_addr_muxed_3_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_6_reg;
  assign c_addr_muxed_3_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_7_reg;
  assign c_addr_muxed_3_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_8_reg;
  assign c_addr_muxed_3_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_9_reg;
  assign c_addr_muxed_3_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_10_reg;
  assign c_addr_muxed_3_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_11_reg;
  assign c_addr_muxed_3_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_12_reg;
  assign c_addr_muxed_3_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_13_reg;
  assign c_addr_muxed_3_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_14_reg;
  assign c_addr_muxed_3_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_3_15_reg;
  assign c_addr_muxed_4_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_0_reg;
  assign c_addr_muxed_4_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_1_reg;
  assign c_addr_muxed_4_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_2_reg;
  assign c_addr_muxed_4_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_3_reg;
  assign c_addr_muxed_4_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_4_reg;
  assign c_addr_muxed_4_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_5_reg;
  assign c_addr_muxed_4_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_6_reg;
  assign c_addr_muxed_4_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_7_reg;
  assign c_addr_muxed_4_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_8_reg;
  assign c_addr_muxed_4_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_9_reg;
  assign c_addr_muxed_4_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_10_reg;
  assign c_addr_muxed_4_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_11_reg;
  assign c_addr_muxed_4_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_12_reg;
  assign c_addr_muxed_4_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_13_reg;
  assign c_addr_muxed_4_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_14_reg;
  assign c_addr_muxed_4_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_4_15_reg;
  assign c_addr_muxed_5_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_0_reg;
  assign c_addr_muxed_5_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_1_reg;
  assign c_addr_muxed_5_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_2_reg;
  assign c_addr_muxed_5_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_3_reg;
  assign c_addr_muxed_5_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_4_reg;
  assign c_addr_muxed_5_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_5_reg;
  assign c_addr_muxed_5_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_6_reg;
  assign c_addr_muxed_5_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_7_reg;
  assign c_addr_muxed_5_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_8_reg;
  assign c_addr_muxed_5_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_9_reg;
  assign c_addr_muxed_5_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_10_reg;
  assign c_addr_muxed_5_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_11_reg;
  assign c_addr_muxed_5_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_12_reg;
  assign c_addr_muxed_5_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_13_reg;
  assign c_addr_muxed_5_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_14_reg;
  assign c_addr_muxed_5_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_5_15_reg;
  assign c_addr_muxed_6_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_0_reg;
  assign c_addr_muxed_6_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_1_reg;
  assign c_addr_muxed_6_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_2_reg;
  assign c_addr_muxed_6_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_3_reg;
  assign c_addr_muxed_6_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_4_reg;
  assign c_addr_muxed_6_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_5_reg;
  assign c_addr_muxed_6_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_6_reg;
  assign c_addr_muxed_6_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_7_reg;
  assign c_addr_muxed_6_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_8_reg;
  assign c_addr_muxed_6_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_9_reg;
  assign c_addr_muxed_6_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_10_reg;
  assign c_addr_muxed_6_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_11_reg;
  assign c_addr_muxed_6_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_12_reg;
  assign c_addr_muxed_6_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_13_reg;
  assign c_addr_muxed_6_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_14_reg;
  assign c_addr_muxed_6_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_6_15_reg;
  assign c_addr_muxed_7_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_0_reg;
  assign c_addr_muxed_7_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_1_reg;
  assign c_addr_muxed_7_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_2_reg;
  assign c_addr_muxed_7_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_3_reg;
  assign c_addr_muxed_7_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_4_reg;
  assign c_addr_muxed_7_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_5_reg;
  assign c_addr_muxed_7_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_6_reg;
  assign c_addr_muxed_7_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_7_reg;
  assign c_addr_muxed_7_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_8_reg;
  assign c_addr_muxed_7_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_9_reg;
  assign c_addr_muxed_7_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_10_reg;
  assign c_addr_muxed_7_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_11_reg;
  assign c_addr_muxed_7_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_12_reg;
  assign c_addr_muxed_7_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_13_reg;
  assign c_addr_muxed_7_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_14_reg;
  assign c_addr_muxed_7_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_7_15_reg;
  assign c_addr_muxed_8_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_0_reg;
  assign c_addr_muxed_8_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_1_reg;
  assign c_addr_muxed_8_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_2_reg;
  assign c_addr_muxed_8_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_3_reg;
  assign c_addr_muxed_8_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_4_reg;
  assign c_addr_muxed_8_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_5_reg;
  assign c_addr_muxed_8_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_6_reg;
  assign c_addr_muxed_8_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_7_reg;
  assign c_addr_muxed_8_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_8_reg;
  assign c_addr_muxed_8_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_9_reg;
  assign c_addr_muxed_8_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_10_reg;
  assign c_addr_muxed_8_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_11_reg;
  assign c_addr_muxed_8_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_12_reg;
  assign c_addr_muxed_8_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_13_reg;
  assign c_addr_muxed_8_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_14_reg;
  assign c_addr_muxed_8_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_8_15_reg;
  assign c_addr_muxed_9_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_0_reg;
  assign c_addr_muxed_9_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_1_reg;
  assign c_addr_muxed_9_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_2_reg;
  assign c_addr_muxed_9_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_3_reg;
  assign c_addr_muxed_9_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_4_reg;
  assign c_addr_muxed_9_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_5_reg;
  assign c_addr_muxed_9_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_6_reg;
  assign c_addr_muxed_9_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_7_reg;
  assign c_addr_muxed_9_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_8_reg;
  assign c_addr_muxed_9_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_9_reg;
  assign c_addr_muxed_9_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_10_reg;
  assign c_addr_muxed_9_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_11_reg;
  assign c_addr_muxed_9_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_12_reg;
  assign c_addr_muxed_9_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_13_reg;
  assign c_addr_muxed_9_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_14_reg;
  assign c_addr_muxed_9_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_9_15_reg;
  assign c_addr_muxed_10_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_0_reg;
  assign c_addr_muxed_10_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_1_reg;
  assign c_addr_muxed_10_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_2_reg;
  assign c_addr_muxed_10_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_3_reg;
  assign c_addr_muxed_10_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_4_reg;
  assign c_addr_muxed_10_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_5_reg;
  assign c_addr_muxed_10_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_6_reg;
  assign c_addr_muxed_10_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_7_reg;
  assign c_addr_muxed_10_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_8_reg;
  assign c_addr_muxed_10_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_9_reg;
  assign c_addr_muxed_10_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_10_reg;
  assign c_addr_muxed_10_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_11_reg;
  assign c_addr_muxed_10_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_12_reg;
  assign c_addr_muxed_10_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_13_reg;
  assign c_addr_muxed_10_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_14_reg;
  assign c_addr_muxed_10_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_10_15_reg;
  assign c_addr_muxed_11_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_0_reg;
  assign c_addr_muxed_11_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_1_reg;
  assign c_addr_muxed_11_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_2_reg;
  assign c_addr_muxed_11_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_3_reg;
  assign c_addr_muxed_11_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_4_reg;
  assign c_addr_muxed_11_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_5_reg;
  assign c_addr_muxed_11_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_6_reg;
  assign c_addr_muxed_11_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_7_reg;
  assign c_addr_muxed_11_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_8_reg;
  assign c_addr_muxed_11_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_9_reg;
  assign c_addr_muxed_11_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_10_reg;
  assign c_addr_muxed_11_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_11_reg;
  assign c_addr_muxed_11_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_12_reg;
  assign c_addr_muxed_11_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_13_reg;
  assign c_addr_muxed_11_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_14_reg;
  assign c_addr_muxed_11_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_11_15_reg;
  assign c_addr_muxed_12_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_0_reg;
  assign c_addr_muxed_12_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_1_reg;
  assign c_addr_muxed_12_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_2_reg;
  assign c_addr_muxed_12_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_3_reg;
  assign c_addr_muxed_12_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_4_reg;
  assign c_addr_muxed_12_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_5_reg;
  assign c_addr_muxed_12_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_6_reg;
  assign c_addr_muxed_12_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_7_reg;
  assign c_addr_muxed_12_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_8_reg;
  assign c_addr_muxed_12_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_9_reg;
  assign c_addr_muxed_12_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_10_reg;
  assign c_addr_muxed_12_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_11_reg;
  assign c_addr_muxed_12_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_12_reg;
  assign c_addr_muxed_12_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_13_reg;
  assign c_addr_muxed_12_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_14_reg;
  assign c_addr_muxed_12_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_12_15_reg;
  assign c_addr_muxed_13_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_0_reg;
  assign c_addr_muxed_13_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_1_reg;
  assign c_addr_muxed_13_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_2_reg;
  assign c_addr_muxed_13_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_3_reg;
  assign c_addr_muxed_13_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_4_reg;
  assign c_addr_muxed_13_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_5_reg;
  assign c_addr_muxed_13_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_6_reg;
  assign c_addr_muxed_13_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_7_reg;
  assign c_addr_muxed_13_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_8_reg;
  assign c_addr_muxed_13_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_9_reg;
  assign c_addr_muxed_13_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_10_reg;
  assign c_addr_muxed_13_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_11_reg;
  assign c_addr_muxed_13_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_12_reg;
  assign c_addr_muxed_13_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_13_reg;
  assign c_addr_muxed_13_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_14_reg;
  assign c_addr_muxed_13_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_13_15_reg;
  assign c_addr_muxed_14_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_0_reg;
  assign c_addr_muxed_14_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_1_reg;
  assign c_addr_muxed_14_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_2_reg;
  assign c_addr_muxed_14_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_3_reg;
  assign c_addr_muxed_14_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_4_reg;
  assign c_addr_muxed_14_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_5_reg;
  assign c_addr_muxed_14_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_6_reg;
  assign c_addr_muxed_14_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_7_reg;
  assign c_addr_muxed_14_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_8_reg;
  assign c_addr_muxed_14_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_9_reg;
  assign c_addr_muxed_14_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_10_reg;
  assign c_addr_muxed_14_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_11_reg;
  assign c_addr_muxed_14_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_12_reg;
  assign c_addr_muxed_14_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_13_reg;
  assign c_addr_muxed_14_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_14_reg;
  assign c_addr_muxed_14_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_14_15_reg;
  assign c_addr_muxed_15_0 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_0_reg;
  assign c_addr_muxed_15_1 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_1_reg;
  assign c_addr_muxed_15_2 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_2_reg;
  assign c_addr_muxed_15_3 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_3_reg;
  assign c_addr_muxed_15_4 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_4_reg;
  assign c_addr_muxed_15_5 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_5_reg;
  assign c_addr_muxed_15_6 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_6_reg;
  assign c_addr_muxed_15_7 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_7_reg;
  assign c_addr_muxed_15_8 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_8_reg;
  assign c_addr_muxed_15_9 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_9_reg;
  assign c_addr_muxed_15_10 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_10_reg;
  assign c_addr_muxed_15_11 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_11_reg;
  assign c_addr_muxed_15_12 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_12_reg;
  assign c_addr_muxed_15_13 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_13_reg;
  assign c_addr_muxed_15_14 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_14_reg;
  assign c_addr_muxed_15_15 = (enable_reading_from_mem) ? addr_pi_reg : c_addr_15_15_reg;

  always @(posedge clk) begin
    if (reset) begin
      c_addr_0_0_reg <= 0;
      c_addr_0_1_reg <= 0;
      c_addr_0_2_reg <= 0;
      c_addr_0_3_reg <= 0;
      c_addr_0_4_reg <= 0;
      c_addr_0_5_reg <= 0;
      c_addr_0_6_reg <= 0;
      c_addr_0_7_reg <= 0;
      c_addr_0_8_reg <= 0;
      c_addr_0_9_reg <= 0;
      c_addr_0_10_reg <= 0;
      c_addr_0_11_reg <= 0;
      c_addr_0_12_reg <= 0;
      c_addr_0_13_reg <= 0;
      c_addr_0_14_reg <= 0;
      c_addr_0_15_reg <= 0;
      c_addr_1_0_reg <= 0;
      c_addr_1_1_reg <= 0;
      c_addr_1_2_reg <= 0;
      c_addr_1_3_reg <= 0;
      c_addr_1_4_reg <= 0;
      c_addr_1_5_reg <= 0;
      c_addr_1_6_reg <= 0;
      c_addr_1_7_reg <= 0;
      c_addr_1_8_reg <= 0;
      c_addr_1_9_reg <= 0;
      c_addr_1_10_reg <= 0;
      c_addr_1_11_reg <= 0;
      c_addr_1_12_reg <= 0;
      c_addr_1_13_reg <= 0;
      c_addr_1_14_reg <= 0;
      c_addr_1_15_reg <= 0;
      c_addr_2_0_reg <= 0;
      c_addr_2_1_reg <= 0;
      c_addr_2_2_reg <= 0;
      c_addr_2_3_reg <= 0;
      c_addr_2_4_reg <= 0;
      c_addr_2_5_reg <= 0;
      c_addr_2_6_reg <= 0;
      c_addr_2_7_reg <= 0;
      c_addr_2_8_reg <= 0;
      c_addr_2_9_reg <= 0;
      c_addr_2_10_reg <= 0;
      c_addr_2_11_reg <= 0;
      c_addr_2_12_reg <= 0;
      c_addr_2_13_reg <= 0;
      c_addr_2_14_reg <= 0;
      c_addr_2_15_reg <= 0;
      c_addr_3_0_reg <= 0;
      c_addr_3_1_reg <= 0;
      c_addr_3_2_reg <= 0;
      c_addr_3_3_reg <= 0;
      c_addr_3_4_reg <= 0;
      c_addr_3_5_reg <= 0;
      c_addr_3_6_reg <= 0;
      c_addr_3_7_reg <= 0;
      c_addr_3_8_reg <= 0;
      c_addr_3_9_reg <= 0;
      c_addr_3_10_reg <= 0;
      c_addr_3_11_reg <= 0;
      c_addr_3_12_reg <= 0;
      c_addr_3_13_reg <= 0;
      c_addr_3_14_reg <= 0;
      c_addr_3_15_reg <= 0;
      c_addr_4_0_reg <= 0;
      c_addr_4_1_reg <= 0;
      c_addr_4_2_reg <= 0;
      c_addr_4_3_reg <= 0;
      c_addr_4_4_reg <= 0;
      c_addr_4_5_reg <= 0;
      c_addr_4_6_reg <= 0;
      c_addr_4_7_reg <= 0;
      c_addr_4_8_reg <= 0;
      c_addr_4_9_reg <= 0;
      c_addr_4_10_reg <= 0;
      c_addr_4_11_reg <= 0;
      c_addr_4_12_reg <= 0;
      c_addr_4_13_reg <= 0;
      c_addr_4_14_reg <= 0;
      c_addr_4_15_reg <= 0;
      c_addr_5_0_reg <= 0;
      c_addr_5_1_reg <= 0;
      c_addr_5_2_reg <= 0;
      c_addr_5_3_reg <= 0;
      c_addr_5_4_reg <= 0;
      c_addr_5_5_reg <= 0;
      c_addr_5_6_reg <= 0;
      c_addr_5_7_reg <= 0;
      c_addr_5_8_reg <= 0;
      c_addr_5_9_reg <= 0;
      c_addr_5_10_reg <= 0;
      c_addr_5_11_reg <= 0;
      c_addr_5_12_reg <= 0;
      c_addr_5_13_reg <= 0;
      c_addr_5_14_reg <= 0;
      c_addr_5_15_reg <= 0;
      c_addr_6_0_reg <= 0;
      c_addr_6_1_reg <= 0;
      c_addr_6_2_reg <= 0;
      c_addr_6_3_reg <= 0;
      c_addr_6_4_reg <= 0;
      c_addr_6_5_reg <= 0;
      c_addr_6_6_reg <= 0;
      c_addr_6_7_reg <= 0;
      c_addr_6_8_reg <= 0;
      c_addr_6_9_reg <= 0;
      c_addr_6_10_reg <= 0;
      c_addr_6_11_reg <= 0;
      c_addr_6_12_reg <= 0;
      c_addr_6_13_reg <= 0;
      c_addr_6_14_reg <= 0;
      c_addr_6_15_reg <= 0;
      c_addr_7_0_reg <= 0;
      c_addr_7_1_reg <= 0;
      c_addr_7_2_reg <= 0;
      c_addr_7_3_reg <= 0;
      c_addr_7_4_reg <= 0;
      c_addr_7_5_reg <= 0;
      c_addr_7_6_reg <= 0;
      c_addr_7_7_reg <= 0;
      c_addr_7_8_reg <= 0;
      c_addr_7_9_reg <= 0;
      c_addr_7_10_reg <= 0;
      c_addr_7_11_reg <= 0;
      c_addr_7_12_reg <= 0;
      c_addr_7_13_reg <= 0;
      c_addr_7_14_reg <= 0;
      c_addr_7_15_reg <= 0;
      c_addr_8_0_reg <= 0;
      c_addr_8_1_reg <= 0;
      c_addr_8_2_reg <= 0;
      c_addr_8_3_reg <= 0;
      c_addr_8_4_reg <= 0;
      c_addr_8_5_reg <= 0;
      c_addr_8_6_reg <= 0;
      c_addr_8_7_reg <= 0;
      c_addr_8_8_reg <= 0;
      c_addr_8_9_reg <= 0;
      c_addr_8_10_reg <= 0;
      c_addr_8_11_reg <= 0;
      c_addr_8_12_reg <= 0;
      c_addr_8_13_reg <= 0;
      c_addr_8_14_reg <= 0;
      c_addr_8_15_reg <= 0;
      c_addr_9_0_reg <= 0;
      c_addr_9_1_reg <= 0;
      c_addr_9_2_reg <= 0;
      c_addr_9_3_reg <= 0;
      c_addr_9_4_reg <= 0;
      c_addr_9_5_reg <= 0;
      c_addr_9_6_reg <= 0;
      c_addr_9_7_reg <= 0;
      c_addr_9_8_reg <= 0;
      c_addr_9_9_reg <= 0;
      c_addr_9_10_reg <= 0;
      c_addr_9_11_reg <= 0;
      c_addr_9_12_reg <= 0;
      c_addr_9_13_reg <= 0;
      c_addr_9_14_reg <= 0;
      c_addr_9_15_reg <= 0;
      c_addr_10_0_reg <= 0;
      c_addr_10_1_reg <= 0;
      c_addr_10_2_reg <= 0;
      c_addr_10_3_reg <= 0;
      c_addr_10_4_reg <= 0;
      c_addr_10_5_reg <= 0;
      c_addr_10_6_reg <= 0;
      c_addr_10_7_reg <= 0;
      c_addr_10_8_reg <= 0;
      c_addr_10_9_reg <= 0;
      c_addr_10_10_reg <= 0;
      c_addr_10_11_reg <= 0;
      c_addr_10_12_reg <= 0;
      c_addr_10_13_reg <= 0;
      c_addr_10_14_reg <= 0;
      c_addr_10_15_reg <= 0;
      c_addr_11_0_reg <= 0;
      c_addr_11_1_reg <= 0;
      c_addr_11_2_reg <= 0;
      c_addr_11_3_reg <= 0;
      c_addr_11_4_reg <= 0;
      c_addr_11_5_reg <= 0;
      c_addr_11_6_reg <= 0;
      c_addr_11_7_reg <= 0;
      c_addr_11_8_reg <= 0;
      c_addr_11_9_reg <= 0;
      c_addr_11_10_reg <= 0;
      c_addr_11_11_reg <= 0;
      c_addr_11_12_reg <= 0;
      c_addr_11_13_reg <= 0;
      c_addr_11_14_reg <= 0;
      c_addr_11_15_reg <= 0;
      c_addr_12_0_reg <= 0;
      c_addr_12_1_reg <= 0;
      c_addr_12_2_reg <= 0;
      c_addr_12_3_reg <= 0;
      c_addr_12_4_reg <= 0;
      c_addr_12_5_reg <= 0;
      c_addr_12_6_reg <= 0;
      c_addr_12_7_reg <= 0;
      c_addr_12_8_reg <= 0;
      c_addr_12_9_reg <= 0;
      c_addr_12_10_reg <= 0;
      c_addr_12_11_reg <= 0;
      c_addr_12_12_reg <= 0;
      c_addr_12_13_reg <= 0;
      c_addr_12_14_reg <= 0;
      c_addr_12_15_reg <= 0;
      c_addr_13_0_reg <= 0;
      c_addr_13_1_reg <= 0;
      c_addr_13_2_reg <= 0;
      c_addr_13_3_reg <= 0;
      c_addr_13_4_reg <= 0;
      c_addr_13_5_reg <= 0;
      c_addr_13_6_reg <= 0;
      c_addr_13_7_reg <= 0;
      c_addr_13_8_reg <= 0;
      c_addr_13_9_reg <= 0;
      c_addr_13_10_reg <= 0;
      c_addr_13_11_reg <= 0;
      c_addr_13_12_reg <= 0;
      c_addr_13_13_reg <= 0;
      c_addr_13_14_reg <= 0;
      c_addr_13_15_reg <= 0;
      c_addr_14_0_reg <= 0;
      c_addr_14_1_reg <= 0;
      c_addr_14_2_reg <= 0;
      c_addr_14_3_reg <= 0;
      c_addr_14_4_reg <= 0;
      c_addr_14_5_reg <= 0;
      c_addr_14_6_reg <= 0;
      c_addr_14_7_reg <= 0;
      c_addr_14_8_reg <= 0;
      c_addr_14_9_reg <= 0;
      c_addr_14_10_reg <= 0;
      c_addr_14_11_reg <= 0;
      c_addr_14_12_reg <= 0;
      c_addr_14_13_reg <= 0;
      c_addr_14_14_reg <= 0;
      c_addr_14_15_reg <= 0;
      c_addr_15_0_reg <= 0;
      c_addr_15_1_reg <= 0;
      c_addr_15_2_reg <= 0;
      c_addr_15_3_reg <= 0;
      c_addr_15_4_reg <= 0;
      c_addr_15_5_reg <= 0;
      c_addr_15_6_reg <= 0;
      c_addr_15_7_reg <= 0;
      c_addr_15_8_reg <= 0;
      c_addr_15_9_reg <= 0;
      c_addr_15_10_reg <= 0;
      c_addr_15_11_reg <= 0;
      c_addr_15_12_reg <= 0;
      c_addr_15_13_reg <= 0;
      c_addr_15_14_reg <= 0;
      c_addr_15_15_reg <= 0;
      c_addr_muxed_0_0_reg <= 0;
      c_addr_muxed_0_1_reg <= 0;
      c_addr_muxed_0_2_reg <= 0;
      c_addr_muxed_0_3_reg <= 0;
      c_addr_muxed_0_4_reg <= 0;
      c_addr_muxed_0_5_reg <= 0;
      c_addr_muxed_0_6_reg <= 0;
      c_addr_muxed_0_7_reg <= 0;
      c_addr_muxed_0_8_reg <= 0;
      c_addr_muxed_0_9_reg <= 0;
      c_addr_muxed_0_10_reg <= 0;
      c_addr_muxed_0_11_reg <= 0;
      c_addr_muxed_0_12_reg <= 0;
      c_addr_muxed_0_13_reg <= 0;
      c_addr_muxed_0_14_reg <= 0;
      c_addr_muxed_0_15_reg <= 0;
      c_addr_muxed_1_0_reg <= 0;
      c_addr_muxed_1_1_reg <= 0;
      c_addr_muxed_1_2_reg <= 0;
      c_addr_muxed_1_3_reg <= 0;
      c_addr_muxed_1_4_reg <= 0;
      c_addr_muxed_1_5_reg <= 0;
      c_addr_muxed_1_6_reg <= 0;
      c_addr_muxed_1_7_reg <= 0;
      c_addr_muxed_1_8_reg <= 0;
      c_addr_muxed_1_9_reg <= 0;
      c_addr_muxed_1_10_reg <= 0;
      c_addr_muxed_1_11_reg <= 0;
      c_addr_muxed_1_12_reg <= 0;
      c_addr_muxed_1_13_reg <= 0;
      c_addr_muxed_1_14_reg <= 0;
      c_addr_muxed_1_15_reg <= 0;
      c_addr_muxed_2_0_reg <= 0;
      c_addr_muxed_2_1_reg <= 0;
      c_addr_muxed_2_2_reg <= 0;
      c_addr_muxed_2_3_reg <= 0;
      c_addr_muxed_2_4_reg <= 0;
      c_addr_muxed_2_5_reg <= 0;
      c_addr_muxed_2_6_reg <= 0;
      c_addr_muxed_2_7_reg <= 0;
      c_addr_muxed_2_8_reg <= 0;
      c_addr_muxed_2_9_reg <= 0;
      c_addr_muxed_2_10_reg <= 0;
      c_addr_muxed_2_11_reg <= 0;
      c_addr_muxed_2_12_reg <= 0;
      c_addr_muxed_2_13_reg <= 0;
      c_addr_muxed_2_14_reg <= 0;
      c_addr_muxed_2_15_reg <= 0;
      c_addr_muxed_3_0_reg <= 0;
      c_addr_muxed_3_1_reg <= 0;
      c_addr_muxed_3_2_reg <= 0;
      c_addr_muxed_3_3_reg <= 0;
      c_addr_muxed_3_4_reg <= 0;
      c_addr_muxed_3_5_reg <= 0;
      c_addr_muxed_3_6_reg <= 0;
      c_addr_muxed_3_7_reg <= 0;
      c_addr_muxed_3_8_reg <= 0;
      c_addr_muxed_3_9_reg <= 0;
      c_addr_muxed_3_10_reg <= 0;
      c_addr_muxed_3_11_reg <= 0;
      c_addr_muxed_3_12_reg <= 0;
      c_addr_muxed_3_13_reg <= 0;
      c_addr_muxed_3_14_reg <= 0;
      c_addr_muxed_3_15_reg <= 0;
      c_addr_muxed_4_0_reg <= 0;
      c_addr_muxed_4_1_reg <= 0;
      c_addr_muxed_4_2_reg <= 0;
      c_addr_muxed_4_3_reg <= 0;
      c_addr_muxed_4_4_reg <= 0;
      c_addr_muxed_4_5_reg <= 0;
      c_addr_muxed_4_6_reg <= 0;
      c_addr_muxed_4_7_reg <= 0;
      c_addr_muxed_4_8_reg <= 0;
      c_addr_muxed_4_9_reg <= 0;
      c_addr_muxed_4_10_reg <= 0;
      c_addr_muxed_4_11_reg <= 0;
      c_addr_muxed_4_12_reg <= 0;
      c_addr_muxed_4_13_reg <= 0;
      c_addr_muxed_4_14_reg <= 0;
      c_addr_muxed_4_15_reg <= 0;
      c_addr_muxed_5_0_reg <= 0;
      c_addr_muxed_5_1_reg <= 0;
      c_addr_muxed_5_2_reg <= 0;
      c_addr_muxed_5_3_reg <= 0;
      c_addr_muxed_5_4_reg <= 0;
      c_addr_muxed_5_5_reg <= 0;
      c_addr_muxed_5_6_reg <= 0;
      c_addr_muxed_5_7_reg <= 0;
      c_addr_muxed_5_8_reg <= 0;
      c_addr_muxed_5_9_reg <= 0;
      c_addr_muxed_5_10_reg <= 0;
      c_addr_muxed_5_11_reg <= 0;
      c_addr_muxed_5_12_reg <= 0;
      c_addr_muxed_5_13_reg <= 0;
      c_addr_muxed_5_14_reg <= 0;
      c_addr_muxed_5_15_reg <= 0;
      c_addr_muxed_6_0_reg <= 0;
      c_addr_muxed_6_1_reg <= 0;
      c_addr_muxed_6_2_reg <= 0;
      c_addr_muxed_6_3_reg <= 0;
      c_addr_muxed_6_4_reg <= 0;
      c_addr_muxed_6_5_reg <= 0;
      c_addr_muxed_6_6_reg <= 0;
      c_addr_muxed_6_7_reg <= 0;
      c_addr_muxed_6_8_reg <= 0;
      c_addr_muxed_6_9_reg <= 0;
      c_addr_muxed_6_10_reg <= 0;
      c_addr_muxed_6_11_reg <= 0;
      c_addr_muxed_6_12_reg <= 0;
      c_addr_muxed_6_13_reg <= 0;
      c_addr_muxed_6_14_reg <= 0;
      c_addr_muxed_6_15_reg <= 0;
      c_addr_muxed_7_0_reg <= 0;
      c_addr_muxed_7_1_reg <= 0;
      c_addr_muxed_7_2_reg <= 0;
      c_addr_muxed_7_3_reg <= 0;
      c_addr_muxed_7_4_reg <= 0;
      c_addr_muxed_7_5_reg <= 0;
      c_addr_muxed_7_6_reg <= 0;
      c_addr_muxed_7_7_reg <= 0;
      c_addr_muxed_7_8_reg <= 0;
      c_addr_muxed_7_9_reg <= 0;
      c_addr_muxed_7_10_reg <= 0;
      c_addr_muxed_7_11_reg <= 0;
      c_addr_muxed_7_12_reg <= 0;
      c_addr_muxed_7_13_reg <= 0;
      c_addr_muxed_7_14_reg <= 0;
      c_addr_muxed_7_15_reg <= 0;
      c_addr_muxed_8_0_reg <= 0;
      c_addr_muxed_8_1_reg <= 0;
      c_addr_muxed_8_2_reg <= 0;
      c_addr_muxed_8_3_reg <= 0;
      c_addr_muxed_8_4_reg <= 0;
      c_addr_muxed_8_5_reg <= 0;
      c_addr_muxed_8_6_reg <= 0;
      c_addr_muxed_8_7_reg <= 0;
      c_addr_muxed_8_8_reg <= 0;
      c_addr_muxed_8_9_reg <= 0;
      c_addr_muxed_8_10_reg <= 0;
      c_addr_muxed_8_11_reg <= 0;
      c_addr_muxed_8_12_reg <= 0;
      c_addr_muxed_8_13_reg <= 0;
      c_addr_muxed_8_14_reg <= 0;
      c_addr_muxed_8_15_reg <= 0;
      c_addr_muxed_9_0_reg <= 0;
      c_addr_muxed_9_1_reg <= 0;
      c_addr_muxed_9_2_reg <= 0;
      c_addr_muxed_9_3_reg <= 0;
      c_addr_muxed_9_4_reg <= 0;
      c_addr_muxed_9_5_reg <= 0;
      c_addr_muxed_9_6_reg <= 0;
      c_addr_muxed_9_7_reg <= 0;
      c_addr_muxed_9_8_reg <= 0;
      c_addr_muxed_9_9_reg <= 0;
      c_addr_muxed_9_10_reg <= 0;
      c_addr_muxed_9_11_reg <= 0;
      c_addr_muxed_9_12_reg <= 0;
      c_addr_muxed_9_13_reg <= 0;
      c_addr_muxed_9_14_reg <= 0;
      c_addr_muxed_9_15_reg <= 0;
      c_addr_muxed_10_0_reg <= 0;
      c_addr_muxed_10_1_reg <= 0;
      c_addr_muxed_10_2_reg <= 0;
      c_addr_muxed_10_3_reg <= 0;
      c_addr_muxed_10_4_reg <= 0;
      c_addr_muxed_10_5_reg <= 0;
      c_addr_muxed_10_6_reg <= 0;
      c_addr_muxed_10_7_reg <= 0;
      c_addr_muxed_10_8_reg <= 0;
      c_addr_muxed_10_9_reg <= 0;
      c_addr_muxed_10_10_reg <= 0;
      c_addr_muxed_10_11_reg <= 0;
      c_addr_muxed_10_12_reg <= 0;
      c_addr_muxed_10_13_reg <= 0;
      c_addr_muxed_10_14_reg <= 0;
      c_addr_muxed_10_15_reg <= 0;
      c_addr_muxed_11_0_reg <= 0;
      c_addr_muxed_11_1_reg <= 0;
      c_addr_muxed_11_2_reg <= 0;
      c_addr_muxed_11_3_reg <= 0;
      c_addr_muxed_11_4_reg <= 0;
      c_addr_muxed_11_5_reg <= 0;
      c_addr_muxed_11_6_reg <= 0;
      c_addr_muxed_11_7_reg <= 0;
      c_addr_muxed_11_8_reg <= 0;
      c_addr_muxed_11_9_reg <= 0;
      c_addr_muxed_11_10_reg <= 0;
      c_addr_muxed_11_11_reg <= 0;
      c_addr_muxed_11_12_reg <= 0;
      c_addr_muxed_11_13_reg <= 0;
      c_addr_muxed_11_14_reg <= 0;
      c_addr_muxed_11_15_reg <= 0;
      c_addr_muxed_12_0_reg <= 0;
      c_addr_muxed_12_1_reg <= 0;
      c_addr_muxed_12_2_reg <= 0;
      c_addr_muxed_12_3_reg <= 0;
      c_addr_muxed_12_4_reg <= 0;
      c_addr_muxed_12_5_reg <= 0;
      c_addr_muxed_12_6_reg <= 0;
      c_addr_muxed_12_7_reg <= 0;
      c_addr_muxed_12_8_reg <= 0;
      c_addr_muxed_12_9_reg <= 0;
      c_addr_muxed_12_10_reg <= 0;
      c_addr_muxed_12_11_reg <= 0;
      c_addr_muxed_12_12_reg <= 0;
      c_addr_muxed_12_13_reg <= 0;
      c_addr_muxed_12_14_reg <= 0;
      c_addr_muxed_12_15_reg <= 0;
      c_addr_muxed_13_0_reg <= 0;
      c_addr_muxed_13_1_reg <= 0;
      c_addr_muxed_13_2_reg <= 0;
      c_addr_muxed_13_3_reg <= 0;
      c_addr_muxed_13_4_reg <= 0;
      c_addr_muxed_13_5_reg <= 0;
      c_addr_muxed_13_6_reg <= 0;
      c_addr_muxed_13_7_reg <= 0;
      c_addr_muxed_13_8_reg <= 0;
      c_addr_muxed_13_9_reg <= 0;
      c_addr_muxed_13_10_reg <= 0;
      c_addr_muxed_13_11_reg <= 0;
      c_addr_muxed_13_12_reg <= 0;
      c_addr_muxed_13_13_reg <= 0;
      c_addr_muxed_13_14_reg <= 0;
      c_addr_muxed_13_15_reg <= 0;
      c_addr_muxed_14_0_reg <= 0;
      c_addr_muxed_14_1_reg <= 0;
      c_addr_muxed_14_2_reg <= 0;
      c_addr_muxed_14_3_reg <= 0;
      c_addr_muxed_14_4_reg <= 0;
      c_addr_muxed_14_5_reg <= 0;
      c_addr_muxed_14_6_reg <= 0;
      c_addr_muxed_14_7_reg <= 0;
      c_addr_muxed_14_8_reg <= 0;
      c_addr_muxed_14_9_reg <= 0;
      c_addr_muxed_14_10_reg <= 0;
      c_addr_muxed_14_11_reg <= 0;
      c_addr_muxed_14_12_reg <= 0;
      c_addr_muxed_14_13_reg <= 0;
      c_addr_muxed_14_14_reg <= 0;
      c_addr_muxed_14_15_reg <= 0;
      c_addr_muxed_15_0_reg <= 0;
      c_addr_muxed_15_1_reg <= 0;
      c_addr_muxed_15_2_reg <= 0;
      c_addr_muxed_15_3_reg <= 0;
      c_addr_muxed_15_4_reg <= 0;
      c_addr_muxed_15_5_reg <= 0;
      c_addr_muxed_15_6_reg <= 0;
      c_addr_muxed_15_7_reg <= 0;
      c_addr_muxed_15_8_reg <= 0;
      c_addr_muxed_15_9_reg <= 0;
      c_addr_muxed_15_10_reg <= 0;
      c_addr_muxed_15_11_reg <= 0;
      c_addr_muxed_15_12_reg <= 0;
      c_addr_muxed_15_13_reg <= 0;
      c_addr_muxed_15_14_reg <= 0;
      c_addr_muxed_15_15_reg <= 0;
    end else begin
      c_addr_0_0_reg <= c_addr_0_0;
      c_addr_0_1_reg <= c_addr_0_1;
      c_addr_0_2_reg <= c_addr_0_2;
      c_addr_0_3_reg <= c_addr_0_3;
      c_addr_0_4_reg <= c_addr_0_4;
      c_addr_0_5_reg <= c_addr_0_5;
      c_addr_0_6_reg <= c_addr_0_6;
      c_addr_0_7_reg <= c_addr_0_7;
      c_addr_0_8_reg <= c_addr_0_8;
      c_addr_0_9_reg <= c_addr_0_9;
      c_addr_0_10_reg <= c_addr_0_10;
      c_addr_0_11_reg <= c_addr_0_11;
      c_addr_0_12_reg <= c_addr_0_12;
      c_addr_0_13_reg <= c_addr_0_13;
      c_addr_0_14_reg <= c_addr_0_14;
      c_addr_0_15_reg <= c_addr_0_15;
      c_addr_1_0_reg <= c_addr_1_0;
      c_addr_1_1_reg <= c_addr_1_1;
      c_addr_1_2_reg <= c_addr_1_2;
      c_addr_1_3_reg <= c_addr_1_3;
      c_addr_1_4_reg <= c_addr_1_4;
      c_addr_1_5_reg <= c_addr_1_5;
      c_addr_1_6_reg <= c_addr_1_6;
      c_addr_1_7_reg <= c_addr_1_7;
      c_addr_1_8_reg <= c_addr_1_8;
      c_addr_1_9_reg <= c_addr_1_9;
      c_addr_1_10_reg <= c_addr_1_10;
      c_addr_1_11_reg <= c_addr_1_11;
      c_addr_1_12_reg <= c_addr_1_12;
      c_addr_1_13_reg <= c_addr_1_13;
      c_addr_1_14_reg <= c_addr_1_14;
      c_addr_1_15_reg <= c_addr_1_15;
      c_addr_2_0_reg <= c_addr_2_0;
      c_addr_2_1_reg <= c_addr_2_1;
      c_addr_2_2_reg <= c_addr_2_2;
      c_addr_2_3_reg <= c_addr_2_3;
      c_addr_2_4_reg <= c_addr_2_4;
      c_addr_2_5_reg <= c_addr_2_5;
      c_addr_2_6_reg <= c_addr_2_6;
      c_addr_2_7_reg <= c_addr_2_7;
      c_addr_2_8_reg <= c_addr_2_8;
      c_addr_2_9_reg <= c_addr_2_9;
      c_addr_2_10_reg <= c_addr_2_10;
      c_addr_2_11_reg <= c_addr_2_11;
      c_addr_2_12_reg <= c_addr_2_12;
      c_addr_2_13_reg <= c_addr_2_13;
      c_addr_2_14_reg <= c_addr_2_14;
      c_addr_2_15_reg <= c_addr_2_15;
      c_addr_3_0_reg <= c_addr_3_0;
      c_addr_3_1_reg <= c_addr_3_1;
      c_addr_3_2_reg <= c_addr_3_2;
      c_addr_3_3_reg <= c_addr_3_3;
      c_addr_3_4_reg <= c_addr_3_4;
      c_addr_3_5_reg <= c_addr_3_5;
      c_addr_3_6_reg <= c_addr_3_6;
      c_addr_3_7_reg <= c_addr_3_7;
      c_addr_3_8_reg <= c_addr_3_8;
      c_addr_3_9_reg <= c_addr_3_9;
      c_addr_3_10_reg <= c_addr_3_10;
      c_addr_3_11_reg <= c_addr_3_11;
      c_addr_3_12_reg <= c_addr_3_12;
      c_addr_3_13_reg <= c_addr_3_13;
      c_addr_3_14_reg <= c_addr_3_14;
      c_addr_3_15_reg <= c_addr_3_15;
      c_addr_4_0_reg <= c_addr_4_0;
      c_addr_4_1_reg <= c_addr_4_1;
      c_addr_4_2_reg <= c_addr_4_2;
      c_addr_4_3_reg <= c_addr_4_3;
      c_addr_4_4_reg <= c_addr_4_4;
      c_addr_4_5_reg <= c_addr_4_5;
      c_addr_4_6_reg <= c_addr_4_6;
      c_addr_4_7_reg <= c_addr_4_7;
      c_addr_4_8_reg <= c_addr_4_8;
      c_addr_4_9_reg <= c_addr_4_9;
      c_addr_4_10_reg <= c_addr_4_10;
      c_addr_4_11_reg <= c_addr_4_11;
      c_addr_4_12_reg <= c_addr_4_12;
      c_addr_4_13_reg <= c_addr_4_13;
      c_addr_4_14_reg <= c_addr_4_14;
      c_addr_4_15_reg <= c_addr_4_15;
      c_addr_5_0_reg <= c_addr_5_0;
      c_addr_5_1_reg <= c_addr_5_1;
      c_addr_5_2_reg <= c_addr_5_2;
      c_addr_5_3_reg <= c_addr_5_3;
      c_addr_5_4_reg <= c_addr_5_4;
      c_addr_5_5_reg <= c_addr_5_5;
      c_addr_5_6_reg <= c_addr_5_6;
      c_addr_5_7_reg <= c_addr_5_7;
      c_addr_5_8_reg <= c_addr_5_8;
      c_addr_5_9_reg <= c_addr_5_9;
      c_addr_5_10_reg <= c_addr_5_10;
      c_addr_5_11_reg <= c_addr_5_11;
      c_addr_5_12_reg <= c_addr_5_12;
      c_addr_5_13_reg <= c_addr_5_13;
      c_addr_5_14_reg <= c_addr_5_14;
      c_addr_5_15_reg <= c_addr_5_15;
      c_addr_6_0_reg <= c_addr_6_0;
      c_addr_6_1_reg <= c_addr_6_1;
      c_addr_6_2_reg <= c_addr_6_2;
      c_addr_6_3_reg <= c_addr_6_3;
      c_addr_6_4_reg <= c_addr_6_4;
      c_addr_6_5_reg <= c_addr_6_5;
      c_addr_6_6_reg <= c_addr_6_6;
      c_addr_6_7_reg <= c_addr_6_7;
      c_addr_6_8_reg <= c_addr_6_8;
      c_addr_6_9_reg <= c_addr_6_9;
      c_addr_6_10_reg <= c_addr_6_10;
      c_addr_6_11_reg <= c_addr_6_11;
      c_addr_6_12_reg <= c_addr_6_12;
      c_addr_6_13_reg <= c_addr_6_13;
      c_addr_6_14_reg <= c_addr_6_14;
      c_addr_6_15_reg <= c_addr_6_15;
      c_addr_7_0_reg <= c_addr_7_0;
      c_addr_7_1_reg <= c_addr_7_1;
      c_addr_7_2_reg <= c_addr_7_2;
      c_addr_7_3_reg <= c_addr_7_3;
      c_addr_7_4_reg <= c_addr_7_4;
      c_addr_7_5_reg <= c_addr_7_5;
      c_addr_7_6_reg <= c_addr_7_6;
      c_addr_7_7_reg <= c_addr_7_7;
      c_addr_7_8_reg <= c_addr_7_8;
      c_addr_7_9_reg <= c_addr_7_9;
      c_addr_7_10_reg <= c_addr_7_10;
      c_addr_7_11_reg <= c_addr_7_11;
      c_addr_7_12_reg <= c_addr_7_12;
      c_addr_7_13_reg <= c_addr_7_13;
      c_addr_7_14_reg <= c_addr_7_14;
      c_addr_7_15_reg <= c_addr_7_15;
      c_addr_8_0_reg <= c_addr_8_0;
      c_addr_8_1_reg <= c_addr_8_1;
      c_addr_8_2_reg <= c_addr_8_2;
      c_addr_8_3_reg <= c_addr_8_3;
      c_addr_8_4_reg <= c_addr_8_4;
      c_addr_8_5_reg <= c_addr_8_5;
      c_addr_8_6_reg <= c_addr_8_6;
      c_addr_8_7_reg <= c_addr_8_7;
      c_addr_8_8_reg <= c_addr_8_8;
      c_addr_8_9_reg <= c_addr_8_9;
      c_addr_8_10_reg <= c_addr_8_10;
      c_addr_8_11_reg <= c_addr_8_11;
      c_addr_8_12_reg <= c_addr_8_12;
      c_addr_8_13_reg <= c_addr_8_13;
      c_addr_8_14_reg <= c_addr_8_14;
      c_addr_8_15_reg <= c_addr_8_15;
      c_addr_9_0_reg <= c_addr_9_0;
      c_addr_9_1_reg <= c_addr_9_1;
      c_addr_9_2_reg <= c_addr_9_2;
      c_addr_9_3_reg <= c_addr_9_3;
      c_addr_9_4_reg <= c_addr_9_4;
      c_addr_9_5_reg <= c_addr_9_5;
      c_addr_9_6_reg <= c_addr_9_6;
      c_addr_9_7_reg <= c_addr_9_7;
      c_addr_9_8_reg <= c_addr_9_8;
      c_addr_9_9_reg <= c_addr_9_9;
      c_addr_9_10_reg <= c_addr_9_10;
      c_addr_9_11_reg <= c_addr_9_11;
      c_addr_9_12_reg <= c_addr_9_12;
      c_addr_9_13_reg <= c_addr_9_13;
      c_addr_9_14_reg <= c_addr_9_14;
      c_addr_9_15_reg <= c_addr_9_15;
      c_addr_10_0_reg <= c_addr_10_0;
      c_addr_10_1_reg <= c_addr_10_1;
      c_addr_10_2_reg <= c_addr_10_2;
      c_addr_10_3_reg <= c_addr_10_3;
      c_addr_10_4_reg <= c_addr_10_4;
      c_addr_10_5_reg <= c_addr_10_5;
      c_addr_10_6_reg <= c_addr_10_6;
      c_addr_10_7_reg <= c_addr_10_7;
      c_addr_10_8_reg <= c_addr_10_8;
      c_addr_10_9_reg <= c_addr_10_9;
      c_addr_10_10_reg <= c_addr_10_10;
      c_addr_10_11_reg <= c_addr_10_11;
      c_addr_10_12_reg <= c_addr_10_12;
      c_addr_10_13_reg <= c_addr_10_13;
      c_addr_10_14_reg <= c_addr_10_14;
      c_addr_10_15_reg <= c_addr_10_15;
      c_addr_11_0_reg <= c_addr_11_0;
      c_addr_11_1_reg <= c_addr_11_1;
      c_addr_11_2_reg <= c_addr_11_2;
      c_addr_11_3_reg <= c_addr_11_3;
      c_addr_11_4_reg <= c_addr_11_4;
      c_addr_11_5_reg <= c_addr_11_5;
      c_addr_11_6_reg <= c_addr_11_6;
      c_addr_11_7_reg <= c_addr_11_7;
      c_addr_11_8_reg <= c_addr_11_8;
      c_addr_11_9_reg <= c_addr_11_9;
      c_addr_11_10_reg <= c_addr_11_10;
      c_addr_11_11_reg <= c_addr_11_11;
      c_addr_11_12_reg <= c_addr_11_12;
      c_addr_11_13_reg <= c_addr_11_13;
      c_addr_11_14_reg <= c_addr_11_14;
      c_addr_11_15_reg <= c_addr_11_15;
      c_addr_12_0_reg <= c_addr_12_0;
      c_addr_12_1_reg <= c_addr_12_1;
      c_addr_12_2_reg <= c_addr_12_2;
      c_addr_12_3_reg <= c_addr_12_3;
      c_addr_12_4_reg <= c_addr_12_4;
      c_addr_12_5_reg <= c_addr_12_5;
      c_addr_12_6_reg <= c_addr_12_6;
      c_addr_12_7_reg <= c_addr_12_7;
      c_addr_12_8_reg <= c_addr_12_8;
      c_addr_12_9_reg <= c_addr_12_9;
      c_addr_12_10_reg <= c_addr_12_10;
      c_addr_12_11_reg <= c_addr_12_11;
      c_addr_12_12_reg <= c_addr_12_12;
      c_addr_12_13_reg <= c_addr_12_13;
      c_addr_12_14_reg <= c_addr_12_14;
      c_addr_12_15_reg <= c_addr_12_15;
      c_addr_13_0_reg <= c_addr_13_0;
      c_addr_13_1_reg <= c_addr_13_1;
      c_addr_13_2_reg <= c_addr_13_2;
      c_addr_13_3_reg <= c_addr_13_3;
      c_addr_13_4_reg <= c_addr_13_4;
      c_addr_13_5_reg <= c_addr_13_5;
      c_addr_13_6_reg <= c_addr_13_6;
      c_addr_13_7_reg <= c_addr_13_7;
      c_addr_13_8_reg <= c_addr_13_8;
      c_addr_13_9_reg <= c_addr_13_9;
      c_addr_13_10_reg <= c_addr_13_10;
      c_addr_13_11_reg <= c_addr_13_11;
      c_addr_13_12_reg <= c_addr_13_12;
      c_addr_13_13_reg <= c_addr_13_13;
      c_addr_13_14_reg <= c_addr_13_14;
      c_addr_13_15_reg <= c_addr_13_15;
      c_addr_14_0_reg <= c_addr_14_0;
      c_addr_14_1_reg <= c_addr_14_1;
      c_addr_14_2_reg <= c_addr_14_2;
      c_addr_14_3_reg <= c_addr_14_3;
      c_addr_14_4_reg <= c_addr_14_4;
      c_addr_14_5_reg <= c_addr_14_5;
      c_addr_14_6_reg <= c_addr_14_6;
      c_addr_14_7_reg <= c_addr_14_7;
      c_addr_14_8_reg <= c_addr_14_8;
      c_addr_14_9_reg <= c_addr_14_9;
      c_addr_14_10_reg <= c_addr_14_10;
      c_addr_14_11_reg <= c_addr_14_11;
      c_addr_14_12_reg <= c_addr_14_12;
      c_addr_14_13_reg <= c_addr_14_13;
      c_addr_14_14_reg <= c_addr_14_14;
      c_addr_14_15_reg <= c_addr_14_15;
      c_addr_15_0_reg <= c_addr_15_0;
      c_addr_15_1_reg <= c_addr_15_1;
      c_addr_15_2_reg <= c_addr_15_2;
      c_addr_15_3_reg <= c_addr_15_3;
      c_addr_15_4_reg <= c_addr_15_4;
      c_addr_15_5_reg <= c_addr_15_5;
      c_addr_15_6_reg <= c_addr_15_6;
      c_addr_15_7_reg <= c_addr_15_7;
      c_addr_15_8_reg <= c_addr_15_8;
      c_addr_15_9_reg <= c_addr_15_9;
      c_addr_15_10_reg <= c_addr_15_10;
      c_addr_15_11_reg <= c_addr_15_11;
      c_addr_15_12_reg <= c_addr_15_12;
      c_addr_15_13_reg <= c_addr_15_13;
      c_addr_15_14_reg <= c_addr_15_14;
      c_addr_15_15_reg <= c_addr_15_15;
      c_addr_muxed_0_0_reg <= c_addr_muxed_0_0;
      c_addr_muxed_0_1_reg <= c_addr_muxed_0_1;
      c_addr_muxed_0_2_reg <= c_addr_muxed_0_2;
      c_addr_muxed_0_3_reg <= c_addr_muxed_0_3;
      c_addr_muxed_0_4_reg <= c_addr_muxed_0_4;
      c_addr_muxed_0_5_reg <= c_addr_muxed_0_5;
      c_addr_muxed_0_6_reg <= c_addr_muxed_0_6;
      c_addr_muxed_0_7_reg <= c_addr_muxed_0_7;
      c_addr_muxed_0_8_reg <= c_addr_muxed_0_8;
      c_addr_muxed_0_9_reg <= c_addr_muxed_0_9;
      c_addr_muxed_0_10_reg <= c_addr_muxed_0_10;
      c_addr_muxed_0_11_reg <= c_addr_muxed_0_11;
      c_addr_muxed_0_12_reg <= c_addr_muxed_0_12;
      c_addr_muxed_0_13_reg <= c_addr_muxed_0_13;
      c_addr_muxed_0_14_reg <= c_addr_muxed_0_14;
      c_addr_muxed_0_15_reg <= c_addr_muxed_0_15;
      c_addr_muxed_1_0_reg <= c_addr_muxed_1_0;
      c_addr_muxed_1_1_reg <= c_addr_muxed_1_1;
      c_addr_muxed_1_2_reg <= c_addr_muxed_1_2;
      c_addr_muxed_1_3_reg <= c_addr_muxed_1_3;
      c_addr_muxed_1_4_reg <= c_addr_muxed_1_4;
      c_addr_muxed_1_5_reg <= c_addr_muxed_1_5;
      c_addr_muxed_1_6_reg <= c_addr_muxed_1_6;
      c_addr_muxed_1_7_reg <= c_addr_muxed_1_7;
      c_addr_muxed_1_8_reg <= c_addr_muxed_1_8;
      c_addr_muxed_1_9_reg <= c_addr_muxed_1_9;
      c_addr_muxed_1_10_reg <= c_addr_muxed_1_10;
      c_addr_muxed_1_11_reg <= c_addr_muxed_1_11;
      c_addr_muxed_1_12_reg <= c_addr_muxed_1_12;
      c_addr_muxed_1_13_reg <= c_addr_muxed_1_13;
      c_addr_muxed_1_14_reg <= c_addr_muxed_1_14;
      c_addr_muxed_1_15_reg <= c_addr_muxed_1_15;
      c_addr_muxed_2_0_reg <= c_addr_muxed_2_0;
      c_addr_muxed_2_1_reg <= c_addr_muxed_2_1;
      c_addr_muxed_2_2_reg <= c_addr_muxed_2_2;
      c_addr_muxed_2_3_reg <= c_addr_muxed_2_3;
      c_addr_muxed_2_4_reg <= c_addr_muxed_2_4;
      c_addr_muxed_2_5_reg <= c_addr_muxed_2_5;
      c_addr_muxed_2_6_reg <= c_addr_muxed_2_6;
      c_addr_muxed_2_7_reg <= c_addr_muxed_2_7;
      c_addr_muxed_2_8_reg <= c_addr_muxed_2_8;
      c_addr_muxed_2_9_reg <= c_addr_muxed_2_9;
      c_addr_muxed_2_10_reg <= c_addr_muxed_2_10;
      c_addr_muxed_2_11_reg <= c_addr_muxed_2_11;
      c_addr_muxed_2_12_reg <= c_addr_muxed_2_12;
      c_addr_muxed_2_13_reg <= c_addr_muxed_2_13;
      c_addr_muxed_2_14_reg <= c_addr_muxed_2_14;
      c_addr_muxed_2_15_reg <= c_addr_muxed_2_15;
      c_addr_muxed_3_0_reg <= c_addr_muxed_3_0;
      c_addr_muxed_3_1_reg <= c_addr_muxed_3_1;
      c_addr_muxed_3_2_reg <= c_addr_muxed_3_2;
      c_addr_muxed_3_3_reg <= c_addr_muxed_3_3;
      c_addr_muxed_3_4_reg <= c_addr_muxed_3_4;
      c_addr_muxed_3_5_reg <= c_addr_muxed_3_5;
      c_addr_muxed_3_6_reg <= c_addr_muxed_3_6;
      c_addr_muxed_3_7_reg <= c_addr_muxed_3_7;
      c_addr_muxed_3_8_reg <= c_addr_muxed_3_8;
      c_addr_muxed_3_9_reg <= c_addr_muxed_3_9;
      c_addr_muxed_3_10_reg <= c_addr_muxed_3_10;
      c_addr_muxed_3_11_reg <= c_addr_muxed_3_11;
      c_addr_muxed_3_12_reg <= c_addr_muxed_3_12;
      c_addr_muxed_3_13_reg <= c_addr_muxed_3_13;
      c_addr_muxed_3_14_reg <= c_addr_muxed_3_14;
      c_addr_muxed_3_15_reg <= c_addr_muxed_3_15;
      c_addr_muxed_4_0_reg <= c_addr_muxed_4_0;
      c_addr_muxed_4_1_reg <= c_addr_muxed_4_1;
      c_addr_muxed_4_2_reg <= c_addr_muxed_4_2;
      c_addr_muxed_4_3_reg <= c_addr_muxed_4_3;
      c_addr_muxed_4_4_reg <= c_addr_muxed_4_4;
      c_addr_muxed_4_5_reg <= c_addr_muxed_4_5;
      c_addr_muxed_4_6_reg <= c_addr_muxed_4_6;
      c_addr_muxed_4_7_reg <= c_addr_muxed_4_7;
      c_addr_muxed_4_8_reg <= c_addr_muxed_4_8;
      c_addr_muxed_4_9_reg <= c_addr_muxed_4_9;
      c_addr_muxed_4_10_reg <= c_addr_muxed_4_10;
      c_addr_muxed_4_11_reg <= c_addr_muxed_4_11;
      c_addr_muxed_4_12_reg <= c_addr_muxed_4_12;
      c_addr_muxed_4_13_reg <= c_addr_muxed_4_13;
      c_addr_muxed_4_14_reg <= c_addr_muxed_4_14;
      c_addr_muxed_4_15_reg <= c_addr_muxed_4_15;
      c_addr_muxed_5_0_reg <= c_addr_muxed_5_0;
      c_addr_muxed_5_1_reg <= c_addr_muxed_5_1;
      c_addr_muxed_5_2_reg <= c_addr_muxed_5_2;
      c_addr_muxed_5_3_reg <= c_addr_muxed_5_3;
      c_addr_muxed_5_4_reg <= c_addr_muxed_5_4;
      c_addr_muxed_5_5_reg <= c_addr_muxed_5_5;
      c_addr_muxed_5_6_reg <= c_addr_muxed_5_6;
      c_addr_muxed_5_7_reg <= c_addr_muxed_5_7;
      c_addr_muxed_5_8_reg <= c_addr_muxed_5_8;
      c_addr_muxed_5_9_reg <= c_addr_muxed_5_9;
      c_addr_muxed_5_10_reg <= c_addr_muxed_5_10;
      c_addr_muxed_5_11_reg <= c_addr_muxed_5_11;
      c_addr_muxed_5_12_reg <= c_addr_muxed_5_12;
      c_addr_muxed_5_13_reg <= c_addr_muxed_5_13;
      c_addr_muxed_5_14_reg <= c_addr_muxed_5_14;
      c_addr_muxed_5_15_reg <= c_addr_muxed_5_15;
      c_addr_muxed_6_0_reg <= c_addr_muxed_6_0;
      c_addr_muxed_6_1_reg <= c_addr_muxed_6_1;
      c_addr_muxed_6_2_reg <= c_addr_muxed_6_2;
      c_addr_muxed_6_3_reg <= c_addr_muxed_6_3;
      c_addr_muxed_6_4_reg <= c_addr_muxed_6_4;
      c_addr_muxed_6_5_reg <= c_addr_muxed_6_5;
      c_addr_muxed_6_6_reg <= c_addr_muxed_6_6;
      c_addr_muxed_6_7_reg <= c_addr_muxed_6_7;
      c_addr_muxed_6_8_reg <= c_addr_muxed_6_8;
      c_addr_muxed_6_9_reg <= c_addr_muxed_6_9;
      c_addr_muxed_6_10_reg <= c_addr_muxed_6_10;
      c_addr_muxed_6_11_reg <= c_addr_muxed_6_11;
      c_addr_muxed_6_12_reg <= c_addr_muxed_6_12;
      c_addr_muxed_6_13_reg <= c_addr_muxed_6_13;
      c_addr_muxed_6_14_reg <= c_addr_muxed_6_14;
      c_addr_muxed_6_15_reg <= c_addr_muxed_6_15;
      c_addr_muxed_7_0_reg <= c_addr_muxed_7_0;
      c_addr_muxed_7_1_reg <= c_addr_muxed_7_1;
      c_addr_muxed_7_2_reg <= c_addr_muxed_7_2;
      c_addr_muxed_7_3_reg <= c_addr_muxed_7_3;
      c_addr_muxed_7_4_reg <= c_addr_muxed_7_4;
      c_addr_muxed_7_5_reg <= c_addr_muxed_7_5;
      c_addr_muxed_7_6_reg <= c_addr_muxed_7_6;
      c_addr_muxed_7_7_reg <= c_addr_muxed_7_7;
      c_addr_muxed_7_8_reg <= c_addr_muxed_7_8;
      c_addr_muxed_7_9_reg <= c_addr_muxed_7_9;
      c_addr_muxed_7_10_reg <= c_addr_muxed_7_10;
      c_addr_muxed_7_11_reg <= c_addr_muxed_7_11;
      c_addr_muxed_7_12_reg <= c_addr_muxed_7_12;
      c_addr_muxed_7_13_reg <= c_addr_muxed_7_13;
      c_addr_muxed_7_14_reg <= c_addr_muxed_7_14;
      c_addr_muxed_7_15_reg <= c_addr_muxed_7_15;
      c_addr_muxed_8_0_reg <= c_addr_muxed_8_0;
      c_addr_muxed_8_1_reg <= c_addr_muxed_8_1;
      c_addr_muxed_8_2_reg <= c_addr_muxed_8_2;
      c_addr_muxed_8_3_reg <= c_addr_muxed_8_3;
      c_addr_muxed_8_4_reg <= c_addr_muxed_8_4;
      c_addr_muxed_8_5_reg <= c_addr_muxed_8_5;
      c_addr_muxed_8_6_reg <= c_addr_muxed_8_6;
      c_addr_muxed_8_7_reg <= c_addr_muxed_8_7;
      c_addr_muxed_8_8_reg <= c_addr_muxed_8_8;
      c_addr_muxed_8_9_reg <= c_addr_muxed_8_9;
      c_addr_muxed_8_10_reg <= c_addr_muxed_8_10;
      c_addr_muxed_8_11_reg <= c_addr_muxed_8_11;
      c_addr_muxed_8_12_reg <= c_addr_muxed_8_12;
      c_addr_muxed_8_13_reg <= c_addr_muxed_8_13;
      c_addr_muxed_8_14_reg <= c_addr_muxed_8_14;
      c_addr_muxed_8_15_reg <= c_addr_muxed_8_15;
      c_addr_muxed_9_0_reg <= c_addr_muxed_9_0;
      c_addr_muxed_9_1_reg <= c_addr_muxed_9_1;
      c_addr_muxed_9_2_reg <= c_addr_muxed_9_2;
      c_addr_muxed_9_3_reg <= c_addr_muxed_9_3;
      c_addr_muxed_9_4_reg <= c_addr_muxed_9_4;
      c_addr_muxed_9_5_reg <= c_addr_muxed_9_5;
      c_addr_muxed_9_6_reg <= c_addr_muxed_9_6;
      c_addr_muxed_9_7_reg <= c_addr_muxed_9_7;
      c_addr_muxed_9_8_reg <= c_addr_muxed_9_8;
      c_addr_muxed_9_9_reg <= c_addr_muxed_9_9;
      c_addr_muxed_9_10_reg <= c_addr_muxed_9_10;
      c_addr_muxed_9_11_reg <= c_addr_muxed_9_11;
      c_addr_muxed_9_12_reg <= c_addr_muxed_9_12;
      c_addr_muxed_9_13_reg <= c_addr_muxed_9_13;
      c_addr_muxed_9_14_reg <= c_addr_muxed_9_14;
      c_addr_muxed_9_15_reg <= c_addr_muxed_9_15;
      c_addr_muxed_10_0_reg <= c_addr_muxed_10_0;
      c_addr_muxed_10_1_reg <= c_addr_muxed_10_1;
      c_addr_muxed_10_2_reg <= c_addr_muxed_10_2;
      c_addr_muxed_10_3_reg <= c_addr_muxed_10_3;
      c_addr_muxed_10_4_reg <= c_addr_muxed_10_4;
      c_addr_muxed_10_5_reg <= c_addr_muxed_10_5;
      c_addr_muxed_10_6_reg <= c_addr_muxed_10_6;
      c_addr_muxed_10_7_reg <= c_addr_muxed_10_7;
      c_addr_muxed_10_8_reg <= c_addr_muxed_10_8;
      c_addr_muxed_10_9_reg <= c_addr_muxed_10_9;
      c_addr_muxed_10_10_reg <= c_addr_muxed_10_10;
      c_addr_muxed_10_11_reg <= c_addr_muxed_10_11;
      c_addr_muxed_10_12_reg <= c_addr_muxed_10_12;
      c_addr_muxed_10_13_reg <= c_addr_muxed_10_13;
      c_addr_muxed_10_14_reg <= c_addr_muxed_10_14;
      c_addr_muxed_10_15_reg <= c_addr_muxed_10_15;
      c_addr_muxed_11_0_reg <= c_addr_muxed_11_0;
      c_addr_muxed_11_1_reg <= c_addr_muxed_11_1;
      c_addr_muxed_11_2_reg <= c_addr_muxed_11_2;
      c_addr_muxed_11_3_reg <= c_addr_muxed_11_3;
      c_addr_muxed_11_4_reg <= c_addr_muxed_11_4;
      c_addr_muxed_11_5_reg <= c_addr_muxed_11_5;
      c_addr_muxed_11_6_reg <= c_addr_muxed_11_6;
      c_addr_muxed_11_7_reg <= c_addr_muxed_11_7;
      c_addr_muxed_11_8_reg <= c_addr_muxed_11_8;
      c_addr_muxed_11_9_reg <= c_addr_muxed_11_9;
      c_addr_muxed_11_10_reg <= c_addr_muxed_11_10;
      c_addr_muxed_11_11_reg <= c_addr_muxed_11_11;
      c_addr_muxed_11_12_reg <= c_addr_muxed_11_12;
      c_addr_muxed_11_13_reg <= c_addr_muxed_11_13;
      c_addr_muxed_11_14_reg <= c_addr_muxed_11_14;
      c_addr_muxed_11_15_reg <= c_addr_muxed_11_15;
      c_addr_muxed_12_0_reg <= c_addr_muxed_12_0;
      c_addr_muxed_12_1_reg <= c_addr_muxed_12_1;
      c_addr_muxed_12_2_reg <= c_addr_muxed_12_2;
      c_addr_muxed_12_3_reg <= c_addr_muxed_12_3;
      c_addr_muxed_12_4_reg <= c_addr_muxed_12_4;
      c_addr_muxed_12_5_reg <= c_addr_muxed_12_5;
      c_addr_muxed_12_6_reg <= c_addr_muxed_12_6;
      c_addr_muxed_12_7_reg <= c_addr_muxed_12_7;
      c_addr_muxed_12_8_reg <= c_addr_muxed_12_8;
      c_addr_muxed_12_9_reg <= c_addr_muxed_12_9;
      c_addr_muxed_12_10_reg <= c_addr_muxed_12_10;
      c_addr_muxed_12_11_reg <= c_addr_muxed_12_11;
      c_addr_muxed_12_12_reg <= c_addr_muxed_12_12;
      c_addr_muxed_12_13_reg <= c_addr_muxed_12_13;
      c_addr_muxed_12_14_reg <= c_addr_muxed_12_14;
      c_addr_muxed_12_15_reg <= c_addr_muxed_12_15;
      c_addr_muxed_13_0_reg <= c_addr_muxed_13_0;
      c_addr_muxed_13_1_reg <= c_addr_muxed_13_1;
      c_addr_muxed_13_2_reg <= c_addr_muxed_13_2;
      c_addr_muxed_13_3_reg <= c_addr_muxed_13_3;
      c_addr_muxed_13_4_reg <= c_addr_muxed_13_4;
      c_addr_muxed_13_5_reg <= c_addr_muxed_13_5;
      c_addr_muxed_13_6_reg <= c_addr_muxed_13_6;
      c_addr_muxed_13_7_reg <= c_addr_muxed_13_7;
      c_addr_muxed_13_8_reg <= c_addr_muxed_13_8;
      c_addr_muxed_13_9_reg <= c_addr_muxed_13_9;
      c_addr_muxed_13_10_reg <= c_addr_muxed_13_10;
      c_addr_muxed_13_11_reg <= c_addr_muxed_13_11;
      c_addr_muxed_13_12_reg <= c_addr_muxed_13_12;
      c_addr_muxed_13_13_reg <= c_addr_muxed_13_13;
      c_addr_muxed_13_14_reg <= c_addr_muxed_13_14;
      c_addr_muxed_13_15_reg <= c_addr_muxed_13_15;
      c_addr_muxed_14_0_reg <= c_addr_muxed_14_0;
      c_addr_muxed_14_1_reg <= c_addr_muxed_14_1;
      c_addr_muxed_14_2_reg <= c_addr_muxed_14_2;
      c_addr_muxed_14_3_reg <= c_addr_muxed_14_3;
      c_addr_muxed_14_4_reg <= c_addr_muxed_14_4;
      c_addr_muxed_14_5_reg <= c_addr_muxed_14_5;
      c_addr_muxed_14_6_reg <= c_addr_muxed_14_6;
      c_addr_muxed_14_7_reg <= c_addr_muxed_14_7;
      c_addr_muxed_14_8_reg <= c_addr_muxed_14_8;
      c_addr_muxed_14_9_reg <= c_addr_muxed_14_9;
      c_addr_muxed_14_10_reg <= c_addr_muxed_14_10;
      c_addr_muxed_14_11_reg <= c_addr_muxed_14_11;
      c_addr_muxed_14_12_reg <= c_addr_muxed_14_12;
      c_addr_muxed_14_13_reg <= c_addr_muxed_14_13;
      c_addr_muxed_14_14_reg <= c_addr_muxed_14_14;
      c_addr_muxed_14_15_reg <= c_addr_muxed_14_15;
      c_addr_muxed_15_0_reg <= c_addr_muxed_15_0;
      c_addr_muxed_15_1_reg <= c_addr_muxed_15_1;
      c_addr_muxed_15_2_reg <= c_addr_muxed_15_2;
      c_addr_muxed_15_3_reg <= c_addr_muxed_15_3;
      c_addr_muxed_15_4_reg <= c_addr_muxed_15_4;
      c_addr_muxed_15_5_reg <= c_addr_muxed_15_5;
      c_addr_muxed_15_6_reg <= c_addr_muxed_15_6;
      c_addr_muxed_15_7_reg <= c_addr_muxed_15_7;
      c_addr_muxed_15_8_reg <= c_addr_muxed_15_8;
      c_addr_muxed_15_9_reg <= c_addr_muxed_15_9;
      c_addr_muxed_15_10_reg <= c_addr_muxed_15_10;
      c_addr_muxed_15_11_reg <= c_addr_muxed_15_11;
      c_addr_muxed_15_12_reg <= c_addr_muxed_15_12;
      c_addr_muxed_15_13_reg <= c_addr_muxed_15_13;
      c_addr_muxed_15_14_reg <= c_addr_muxed_15_14;
      c_addr_muxed_15_15_reg <= c_addr_muxed_15_15;
    end
  end
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_0_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_1_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_2_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_3_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_4_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_5_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_6_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_7_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_8_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_9_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_10_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_11_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_12_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_13_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_14_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat_15_15;

///////////////// ORing the data ///////////////////
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] data_from_out_mat;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_0;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_1;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_2;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_3;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_4;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_5;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_6;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_7;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_8;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_9;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_10;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_11;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_12;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_13;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_14;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_15;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_16;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_17;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_18;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_19;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_20;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_21;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_22;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_23;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_24;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_25;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_26;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_27;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_28;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_29;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_30;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_31;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_32;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_33;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_34;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_35;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_36;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_37;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_38;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_39;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_40;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_41;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_42;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_43;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_44;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_45;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_46;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_47;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_48;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_49;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_50;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_51;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_52;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_53;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_54;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_55;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_56;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_57;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_58;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_59;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_60;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_61;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_62;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_63;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_64;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_65;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_66;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_67;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_68;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_69;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_70;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_71;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_72;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_73;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_74;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_75;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_76;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_77;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_78;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_79;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_80;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_81;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_82;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_83;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_84;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_85;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_86;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_87;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_88;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_89;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_90;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_91;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_92;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_93;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_94;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_95;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_96;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_97;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_98;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_99;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_100;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_101;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_102;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_103;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_104;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_105;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_106;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_107;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_108;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_109;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_110;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_111;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_112;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_113;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_114;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_115;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_116;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_117;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_118;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_119;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_120;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_121;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_122;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_123;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_124;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_125;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_126;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_127;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_128;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_129;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_130;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_131;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_132;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_133;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_134;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_135;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_136;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_137;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_138;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_139;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_140;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_141;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_142;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_143;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_144;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_145;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_146;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_147;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_148;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_149;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_150;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_151;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_152;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_153;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_154;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_155;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_156;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_157;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_158;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_159;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_160;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_161;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_162;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_163;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_164;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_165;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_166;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_167;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_168;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_169;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_170;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_171;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_172;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_173;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_174;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_175;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_176;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_177;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_178;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_179;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_180;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_181;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_182;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_183;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_184;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_185;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_186;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_187;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_188;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_189;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_190;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_191;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_192;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_193;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_194;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_195;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_196;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_197;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_198;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_199;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_200;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_201;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_202;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_203;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_204;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_205;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_206;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_207;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_208;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_209;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_210;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_211;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_212;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_213;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_214;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_215;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_216;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_217;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_218;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_219;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_220;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_221;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_222;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_223;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_224;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_225;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_226;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_227;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_228;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_229;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_230;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_231;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_232;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_233;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_234;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_235;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_236;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_237;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_238;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_239;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_240;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_241;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_242;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_243;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_244;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_245;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_246;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_247;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_248;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_249;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_250;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_251;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_252;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_253;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_254;
  reg [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_reg_255;
  always @(posedge clk) begin
    if (reset) begin
      c_reg_0 <= 0;
      c_reg_1 <= 0;
      c_reg_2 <= 0;
      c_reg_3 <= 0;
      c_reg_4 <= 0;
      c_reg_5 <= 0;
      c_reg_6 <= 0;
      c_reg_7 <= 0;
      c_reg_8 <= 0;
      c_reg_9 <= 0;
      c_reg_10 <= 0;
      c_reg_11 <= 0;
      c_reg_12 <= 0;
      c_reg_13 <= 0;
      c_reg_14 <= 0;
      c_reg_15 <= 0;
      c_reg_16 <= 0;
      c_reg_17 <= 0;
      c_reg_18 <= 0;
      c_reg_19 <= 0;
      c_reg_20 <= 0;
      c_reg_21 <= 0;
      c_reg_22 <= 0;
      c_reg_23 <= 0;
      c_reg_24 <= 0;
      c_reg_25 <= 0;
      c_reg_26 <= 0;
      c_reg_27 <= 0;
      c_reg_28 <= 0;
      c_reg_29 <= 0;
      c_reg_30 <= 0;
      c_reg_31 <= 0;
      c_reg_32 <= 0;
      c_reg_33 <= 0;
      c_reg_34 <= 0;
      c_reg_35 <= 0;
      c_reg_36 <= 0;
      c_reg_37 <= 0;
      c_reg_38 <= 0;
      c_reg_39 <= 0;
      c_reg_40 <= 0;
      c_reg_41 <= 0;
      c_reg_42 <= 0;
      c_reg_43 <= 0;
      c_reg_44 <= 0;
      c_reg_45 <= 0;
      c_reg_46 <= 0;
      c_reg_47 <= 0;
      c_reg_48 <= 0;
      c_reg_49 <= 0;
      c_reg_50 <= 0;
      c_reg_51 <= 0;
      c_reg_52 <= 0;
      c_reg_53 <= 0;
      c_reg_54 <= 0;
      c_reg_55 <= 0;
      c_reg_56 <= 0;
      c_reg_57 <= 0;
      c_reg_58 <= 0;
      c_reg_59 <= 0;
      c_reg_60 <= 0;
      c_reg_61 <= 0;
      c_reg_62 <= 0;
      c_reg_63 <= 0;
      c_reg_64 <= 0;
      c_reg_65 <= 0;
      c_reg_66 <= 0;
      c_reg_67 <= 0;
      c_reg_68 <= 0;
      c_reg_69 <= 0;
      c_reg_70 <= 0;
      c_reg_71 <= 0;
      c_reg_72 <= 0;
      c_reg_73 <= 0;
      c_reg_74 <= 0;
      c_reg_75 <= 0;
      c_reg_76 <= 0;
      c_reg_77 <= 0;
      c_reg_78 <= 0;
      c_reg_79 <= 0;
      c_reg_80 <= 0;
      c_reg_81 <= 0;
      c_reg_82 <= 0;
      c_reg_83 <= 0;
      c_reg_84 <= 0;
      c_reg_85 <= 0;
      c_reg_86 <= 0;
      c_reg_87 <= 0;
      c_reg_88 <= 0;
      c_reg_89 <= 0;
      c_reg_90 <= 0;
      c_reg_91 <= 0;
      c_reg_92 <= 0;
      c_reg_93 <= 0;
      c_reg_94 <= 0;
      c_reg_95 <= 0;
      c_reg_96 <= 0;
      c_reg_97 <= 0;
      c_reg_98 <= 0;
      c_reg_99 <= 0;
      c_reg_100 <= 0;
      c_reg_101 <= 0;
      c_reg_102 <= 0;
      c_reg_103 <= 0;
      c_reg_104 <= 0;
      c_reg_105 <= 0;
      c_reg_106 <= 0;
      c_reg_107 <= 0;
      c_reg_108 <= 0;
      c_reg_109 <= 0;
      c_reg_110 <= 0;
      c_reg_111 <= 0;
      c_reg_112 <= 0;
      c_reg_113 <= 0;
      c_reg_114 <= 0;
      c_reg_115 <= 0;
      c_reg_116 <= 0;
      c_reg_117 <= 0;
      c_reg_118 <= 0;
      c_reg_119 <= 0;
      c_reg_120 <= 0;
      c_reg_121 <= 0;
      c_reg_122 <= 0;
      c_reg_123 <= 0;
      c_reg_124 <= 0;
      c_reg_125 <= 0;
      c_reg_126 <= 0;
      c_reg_127 <= 0;
      c_reg_128 <= 0;
      c_reg_129 <= 0;
      c_reg_130 <= 0;
      c_reg_131 <= 0;
      c_reg_132 <= 0;
      c_reg_133 <= 0;
      c_reg_134 <= 0;
      c_reg_135 <= 0;
      c_reg_136 <= 0;
      c_reg_137 <= 0;
      c_reg_138 <= 0;
      c_reg_139 <= 0;
      c_reg_140 <= 0;
      c_reg_141 <= 0;
      c_reg_142 <= 0;
      c_reg_143 <= 0;
      c_reg_144 <= 0;
      c_reg_145 <= 0;
      c_reg_146 <= 0;
      c_reg_147 <= 0;
      c_reg_148 <= 0;
      c_reg_149 <= 0;
      c_reg_150 <= 0;
      c_reg_151 <= 0;
      c_reg_152 <= 0;
      c_reg_153 <= 0;
      c_reg_154 <= 0;
      c_reg_155 <= 0;
      c_reg_156 <= 0;
      c_reg_157 <= 0;
      c_reg_158 <= 0;
      c_reg_159 <= 0;
      c_reg_160 <= 0;
      c_reg_161 <= 0;
      c_reg_162 <= 0;
      c_reg_163 <= 0;
      c_reg_164 <= 0;
      c_reg_165 <= 0;
      c_reg_166 <= 0;
      c_reg_167 <= 0;
      c_reg_168 <= 0;
      c_reg_169 <= 0;
      c_reg_170 <= 0;
      c_reg_171 <= 0;
      c_reg_172 <= 0;
      c_reg_173 <= 0;
      c_reg_174 <= 0;
      c_reg_175 <= 0;
      c_reg_176 <= 0;
      c_reg_177 <= 0;
      c_reg_178 <= 0;
      c_reg_179 <= 0;
      c_reg_180 <= 0;
      c_reg_181 <= 0;
      c_reg_182 <= 0;
      c_reg_183 <= 0;
      c_reg_184 <= 0;
      c_reg_185 <= 0;
      c_reg_186 <= 0;
      c_reg_187 <= 0;
      c_reg_188 <= 0;
      c_reg_189 <= 0;
      c_reg_190 <= 0;
      c_reg_191 <= 0;
      c_reg_192 <= 0;
      c_reg_193 <= 0;
      c_reg_194 <= 0;
      c_reg_195 <= 0;
      c_reg_196 <= 0;
      c_reg_197 <= 0;
      c_reg_198 <= 0;
      c_reg_199 <= 0;
      c_reg_200 <= 0;
      c_reg_201 <= 0;
      c_reg_202 <= 0;
      c_reg_203 <= 0;
      c_reg_204 <= 0;
      c_reg_205 <= 0;
      c_reg_206 <= 0;
      c_reg_207 <= 0;
      c_reg_208 <= 0;
      c_reg_209 <= 0;
      c_reg_210 <= 0;
      c_reg_211 <= 0;
      c_reg_212 <= 0;
      c_reg_213 <= 0;
      c_reg_214 <= 0;
      c_reg_215 <= 0;
      c_reg_216 <= 0;
      c_reg_217 <= 0;
      c_reg_218 <= 0;
      c_reg_219 <= 0;
      c_reg_220 <= 0;
      c_reg_221 <= 0;
      c_reg_222 <= 0;
      c_reg_223 <= 0;
      c_reg_224 <= 0;
      c_reg_225 <= 0;
      c_reg_226 <= 0;
      c_reg_227 <= 0;
      c_reg_228 <= 0;
      c_reg_229 <= 0;
      c_reg_230 <= 0;
      c_reg_231 <= 0;
      c_reg_232 <= 0;
      c_reg_233 <= 0;
      c_reg_234 <= 0;
      c_reg_235 <= 0;
      c_reg_236 <= 0;
      c_reg_237 <= 0;
      c_reg_238 <= 0;
      c_reg_239 <= 0;
      c_reg_240 <= 0;
      c_reg_241 <= 0;
      c_reg_242 <= 0;
      c_reg_243 <= 0;
      c_reg_244 <= 0;
      c_reg_245 <= 0;
      c_reg_246 <= 0;
      c_reg_247 <= 0;
      c_reg_248 <= 0;
      c_reg_249 <= 0;
      c_reg_250 <= 0;
      c_reg_251 <= 0;
      c_reg_252 <= 0;
      c_reg_253 <= 0;
      c_reg_254 <= 0;
      c_reg_255 <= 0;
    end else begin
      c_reg_0 <= data_from_out_mat_0_0;
      c_reg_1 <= c_reg_0 | data_from_out_mat_0_1;
      c_reg_2 <= c_reg_1 | data_from_out_mat_0_2;
      c_reg_3 <= c_reg_2 | data_from_out_mat_0_3;
      c_reg_4 <= c_reg_3 | data_from_out_mat_0_4;
      c_reg_5 <= c_reg_4 | data_from_out_mat_0_5;
      c_reg_6 <= c_reg_5 | data_from_out_mat_0_6;
      c_reg_7 <= c_reg_6 | data_from_out_mat_0_7;
      c_reg_8 <= c_reg_7 | data_from_out_mat_0_8;
      c_reg_9 <= c_reg_8 | data_from_out_mat_0_9;
      c_reg_10 <= c_reg_9 | data_from_out_mat_0_10;
      c_reg_11 <= c_reg_10 | data_from_out_mat_0_11;
      c_reg_12 <= c_reg_11 | data_from_out_mat_0_12;
      c_reg_13 <= c_reg_12 | data_from_out_mat_0_13;
      c_reg_14 <= c_reg_13 | data_from_out_mat_0_14;
      c_reg_15 <= c_reg_14 | data_from_out_mat_0_15;
      c_reg_16 <= c_reg_15 | data_from_out_mat_1_0;
      c_reg_17 <= c_reg_16 | data_from_out_mat_1_1;
      c_reg_18 <= c_reg_17 | data_from_out_mat_1_2;
      c_reg_19 <= c_reg_18 | data_from_out_mat_1_3;
      c_reg_20 <= c_reg_19 | data_from_out_mat_1_4;
      c_reg_21 <= c_reg_20 | data_from_out_mat_1_5;
      c_reg_22 <= c_reg_21 | data_from_out_mat_1_6;
      c_reg_23 <= c_reg_22 | data_from_out_mat_1_7;
      c_reg_24 <= c_reg_23 | data_from_out_mat_1_8;
      c_reg_25 <= c_reg_24 | data_from_out_mat_1_9;
      c_reg_26 <= c_reg_25 | data_from_out_mat_1_10;
      c_reg_27 <= c_reg_26 | data_from_out_mat_1_11;
      c_reg_28 <= c_reg_27 | data_from_out_mat_1_12;
      c_reg_29 <= c_reg_28 | data_from_out_mat_1_13;
      c_reg_30 <= c_reg_29 | data_from_out_mat_1_14;
      c_reg_31 <= c_reg_30 | data_from_out_mat_1_15;
      c_reg_32 <= c_reg_31 | data_from_out_mat_2_0;
      c_reg_33 <= c_reg_32 | data_from_out_mat_2_1;
      c_reg_34 <= c_reg_33 | data_from_out_mat_2_2;
      c_reg_35 <= c_reg_34 | data_from_out_mat_2_3;
      c_reg_36 <= c_reg_35 | data_from_out_mat_2_4;
      c_reg_37 <= c_reg_36 | data_from_out_mat_2_5;
      c_reg_38 <= c_reg_37 | data_from_out_mat_2_6;
      c_reg_39 <= c_reg_38 | data_from_out_mat_2_7;
      c_reg_40 <= c_reg_39 | data_from_out_mat_2_8;
      c_reg_41 <= c_reg_40 | data_from_out_mat_2_9;
      c_reg_42 <= c_reg_41 | data_from_out_mat_2_10;
      c_reg_43 <= c_reg_42 | data_from_out_mat_2_11;
      c_reg_44 <= c_reg_43 | data_from_out_mat_2_12;
      c_reg_45 <= c_reg_44 | data_from_out_mat_2_13;
      c_reg_46 <= c_reg_45 | data_from_out_mat_2_14;
      c_reg_47 <= c_reg_46 | data_from_out_mat_2_15;
      c_reg_48 <= c_reg_47 | data_from_out_mat_3_0;
      c_reg_49 <= c_reg_48 | data_from_out_mat_3_1;
      c_reg_50 <= c_reg_49 | data_from_out_mat_3_2;
      c_reg_51 <= c_reg_50 | data_from_out_mat_3_3;
      c_reg_52 <= c_reg_51 | data_from_out_mat_3_4;
      c_reg_53 <= c_reg_52 | data_from_out_mat_3_5;
      c_reg_54 <= c_reg_53 | data_from_out_mat_3_6;
      c_reg_55 <= c_reg_54 | data_from_out_mat_3_7;
      c_reg_56 <= c_reg_55 | data_from_out_mat_3_8;
      c_reg_57 <= c_reg_56 | data_from_out_mat_3_9;
      c_reg_58 <= c_reg_57 | data_from_out_mat_3_10;
      c_reg_59 <= c_reg_58 | data_from_out_mat_3_11;
      c_reg_60 <= c_reg_59 | data_from_out_mat_3_12;
      c_reg_61 <= c_reg_60 | data_from_out_mat_3_13;
      c_reg_62 <= c_reg_61 | data_from_out_mat_3_14;
      c_reg_63 <= c_reg_62 | data_from_out_mat_3_15;
      c_reg_64 <= c_reg_63 | data_from_out_mat_4_0;
      c_reg_65 <= c_reg_64 | data_from_out_mat_4_1;
      c_reg_66 <= c_reg_65 | data_from_out_mat_4_2;
      c_reg_67 <= c_reg_66 | data_from_out_mat_4_3;
      c_reg_68 <= c_reg_67 | data_from_out_mat_4_4;
      c_reg_69 <= c_reg_68 | data_from_out_mat_4_5;
      c_reg_70 <= c_reg_69 | data_from_out_mat_4_6;
      c_reg_71 <= c_reg_70 | data_from_out_mat_4_7;
      c_reg_72 <= c_reg_71 | data_from_out_mat_4_8;
      c_reg_73 <= c_reg_72 | data_from_out_mat_4_9;
      c_reg_74 <= c_reg_73 | data_from_out_mat_4_10;
      c_reg_75 <= c_reg_74 | data_from_out_mat_4_11;
      c_reg_76 <= c_reg_75 | data_from_out_mat_4_12;
      c_reg_77 <= c_reg_76 | data_from_out_mat_4_13;
      c_reg_78 <= c_reg_77 | data_from_out_mat_4_14;
      c_reg_79 <= c_reg_78 | data_from_out_mat_4_15;
      c_reg_80 <= c_reg_79 | data_from_out_mat_5_0;
      c_reg_81 <= c_reg_80 | data_from_out_mat_5_1;
      c_reg_82 <= c_reg_81 | data_from_out_mat_5_2;
      c_reg_83 <= c_reg_82 | data_from_out_mat_5_3;
      c_reg_84 <= c_reg_83 | data_from_out_mat_5_4;
      c_reg_85 <= c_reg_84 | data_from_out_mat_5_5;
      c_reg_86 <= c_reg_85 | data_from_out_mat_5_6;
      c_reg_87 <= c_reg_86 | data_from_out_mat_5_7;
      c_reg_88 <= c_reg_87 | data_from_out_mat_5_8;
      c_reg_89 <= c_reg_88 | data_from_out_mat_5_9;
      c_reg_90 <= c_reg_89 | data_from_out_mat_5_10;
      c_reg_91 <= c_reg_90 | data_from_out_mat_5_11;
      c_reg_92 <= c_reg_91 | data_from_out_mat_5_12;
      c_reg_93 <= c_reg_92 | data_from_out_mat_5_13;
      c_reg_94 <= c_reg_93 | data_from_out_mat_5_14;
      c_reg_95 <= c_reg_94 | data_from_out_mat_5_15;
      c_reg_96 <= c_reg_95 | data_from_out_mat_6_0;
      c_reg_97 <= c_reg_96 | data_from_out_mat_6_1;
      c_reg_98 <= c_reg_97 | data_from_out_mat_6_2;
      c_reg_99 <= c_reg_98 | data_from_out_mat_6_3;
      c_reg_100 <= c_reg_99 | data_from_out_mat_6_4;
      c_reg_101 <= c_reg_100 | data_from_out_mat_6_5;
      c_reg_102 <= c_reg_101 | data_from_out_mat_6_6;
      c_reg_103 <= c_reg_102 | data_from_out_mat_6_7;
      c_reg_104 <= c_reg_103 | data_from_out_mat_6_8;
      c_reg_105 <= c_reg_104 | data_from_out_mat_6_9;
      c_reg_106 <= c_reg_105 | data_from_out_mat_6_10;
      c_reg_107 <= c_reg_106 | data_from_out_mat_6_11;
      c_reg_108 <= c_reg_107 | data_from_out_mat_6_12;
      c_reg_109 <= c_reg_108 | data_from_out_mat_6_13;
      c_reg_110 <= c_reg_109 | data_from_out_mat_6_14;
      c_reg_111 <= c_reg_110 | data_from_out_mat_6_15;
      c_reg_112 <= c_reg_111 | data_from_out_mat_7_0;
      c_reg_113 <= c_reg_112 | data_from_out_mat_7_1;
      c_reg_114 <= c_reg_113 | data_from_out_mat_7_2;
      c_reg_115 <= c_reg_114 | data_from_out_mat_7_3;
      c_reg_116 <= c_reg_115 | data_from_out_mat_7_4;
      c_reg_117 <= c_reg_116 | data_from_out_mat_7_5;
      c_reg_118 <= c_reg_117 | data_from_out_mat_7_6;
      c_reg_119 <= c_reg_118 | data_from_out_mat_7_7;
      c_reg_120 <= c_reg_119 | data_from_out_mat_7_8;
      c_reg_121 <= c_reg_120 | data_from_out_mat_7_9;
      c_reg_122 <= c_reg_121 | data_from_out_mat_7_10;
      c_reg_123 <= c_reg_122 | data_from_out_mat_7_11;
      c_reg_124 <= c_reg_123 | data_from_out_mat_7_12;
      c_reg_125 <= c_reg_124 | data_from_out_mat_7_13;
      c_reg_126 <= c_reg_125 | data_from_out_mat_7_14;
      c_reg_127 <= c_reg_126 | data_from_out_mat_7_15;
      c_reg_128 <= c_reg_127 | data_from_out_mat_8_0;
      c_reg_129 <= c_reg_128 | data_from_out_mat_8_1;
      c_reg_130 <= c_reg_129 | data_from_out_mat_8_2;
      c_reg_131 <= c_reg_130 | data_from_out_mat_8_3;
      c_reg_132 <= c_reg_131 | data_from_out_mat_8_4;
      c_reg_133 <= c_reg_132 | data_from_out_mat_8_5;
      c_reg_134 <= c_reg_133 | data_from_out_mat_8_6;
      c_reg_135 <= c_reg_134 | data_from_out_mat_8_7;
      c_reg_136 <= c_reg_135 | data_from_out_mat_8_8;
      c_reg_137 <= c_reg_136 | data_from_out_mat_8_9;
      c_reg_138 <= c_reg_137 | data_from_out_mat_8_10;
      c_reg_139 <= c_reg_138 | data_from_out_mat_8_11;
      c_reg_140 <= c_reg_139 | data_from_out_mat_8_12;
      c_reg_141 <= c_reg_140 | data_from_out_mat_8_13;
      c_reg_142 <= c_reg_141 | data_from_out_mat_8_14;
      c_reg_143 <= c_reg_142 | data_from_out_mat_8_15;
      c_reg_144 <= c_reg_143 | data_from_out_mat_9_0;
      c_reg_145 <= c_reg_144 | data_from_out_mat_9_1;
      c_reg_146 <= c_reg_145 | data_from_out_mat_9_2;
      c_reg_147 <= c_reg_146 | data_from_out_mat_9_3;
      c_reg_148 <= c_reg_147 | data_from_out_mat_9_4;
      c_reg_149 <= c_reg_148 | data_from_out_mat_9_5;
      c_reg_150 <= c_reg_149 | data_from_out_mat_9_6;
      c_reg_151 <= c_reg_150 | data_from_out_mat_9_7;
      c_reg_152 <= c_reg_151 | data_from_out_mat_9_8;
      c_reg_153 <= c_reg_152 | data_from_out_mat_9_9;
      c_reg_154 <= c_reg_153 | data_from_out_mat_9_10;
      c_reg_155 <= c_reg_154 | data_from_out_mat_9_11;
      c_reg_156 <= c_reg_155 | data_from_out_mat_9_12;
      c_reg_157 <= c_reg_156 | data_from_out_mat_9_13;
      c_reg_158 <= c_reg_157 | data_from_out_mat_9_14;
      c_reg_159 <= c_reg_158 | data_from_out_mat_9_15;
      c_reg_160 <= c_reg_159 | data_from_out_mat_10_0;
      c_reg_161 <= c_reg_160 | data_from_out_mat_10_1;
      c_reg_162 <= c_reg_161 | data_from_out_mat_10_2;
      c_reg_163 <= c_reg_162 | data_from_out_mat_10_3;
      c_reg_164 <= c_reg_163 | data_from_out_mat_10_4;
      c_reg_165 <= c_reg_164 | data_from_out_mat_10_5;
      c_reg_166 <= c_reg_165 | data_from_out_mat_10_6;
      c_reg_167 <= c_reg_166 | data_from_out_mat_10_7;
      c_reg_168 <= c_reg_167 | data_from_out_mat_10_8;
      c_reg_169 <= c_reg_168 | data_from_out_mat_10_9;
      c_reg_170 <= c_reg_169 | data_from_out_mat_10_10;
      c_reg_171 <= c_reg_170 | data_from_out_mat_10_11;
      c_reg_172 <= c_reg_171 | data_from_out_mat_10_12;
      c_reg_173 <= c_reg_172 | data_from_out_mat_10_13;
      c_reg_174 <= c_reg_173 | data_from_out_mat_10_14;
      c_reg_175 <= c_reg_174 | data_from_out_mat_10_15;
      c_reg_176 <= c_reg_175 | data_from_out_mat_11_0;
      c_reg_177 <= c_reg_176 | data_from_out_mat_11_1;
      c_reg_178 <= c_reg_177 | data_from_out_mat_11_2;
      c_reg_179 <= c_reg_178 | data_from_out_mat_11_3;
      c_reg_180 <= c_reg_179 | data_from_out_mat_11_4;
      c_reg_181 <= c_reg_180 | data_from_out_mat_11_5;
      c_reg_182 <= c_reg_181 | data_from_out_mat_11_6;
      c_reg_183 <= c_reg_182 | data_from_out_mat_11_7;
      c_reg_184 <= c_reg_183 | data_from_out_mat_11_8;
      c_reg_185 <= c_reg_184 | data_from_out_mat_11_9;
      c_reg_186 <= c_reg_185 | data_from_out_mat_11_10;
      c_reg_187 <= c_reg_186 | data_from_out_mat_11_11;
      c_reg_188 <= c_reg_187 | data_from_out_mat_11_12;
      c_reg_189 <= c_reg_188 | data_from_out_mat_11_13;
      c_reg_190 <= c_reg_189 | data_from_out_mat_11_14;
      c_reg_191 <= c_reg_190 | data_from_out_mat_11_15;
      c_reg_192 <= c_reg_191 | data_from_out_mat_12_0;
      c_reg_193 <= c_reg_192 | data_from_out_mat_12_1;
      c_reg_194 <= c_reg_193 | data_from_out_mat_12_2;
      c_reg_195 <= c_reg_194 | data_from_out_mat_12_3;
      c_reg_196 <= c_reg_195 | data_from_out_mat_12_4;
      c_reg_197 <= c_reg_196 | data_from_out_mat_12_5;
      c_reg_198 <= c_reg_197 | data_from_out_mat_12_6;
      c_reg_199 <= c_reg_198 | data_from_out_mat_12_7;
      c_reg_200 <= c_reg_199 | data_from_out_mat_12_8;
      c_reg_201 <= c_reg_200 | data_from_out_mat_12_9;
      c_reg_202 <= c_reg_201 | data_from_out_mat_12_10;
      c_reg_203 <= c_reg_202 | data_from_out_mat_12_11;
      c_reg_204 <= c_reg_203 | data_from_out_mat_12_12;
      c_reg_205 <= c_reg_204 | data_from_out_mat_12_13;
      c_reg_206 <= c_reg_205 | data_from_out_mat_12_14;
      c_reg_207 <= c_reg_206 | data_from_out_mat_12_15;
      c_reg_208 <= c_reg_207 | data_from_out_mat_13_0;
      c_reg_209 <= c_reg_208 | data_from_out_mat_13_1;
      c_reg_210 <= c_reg_209 | data_from_out_mat_13_2;
      c_reg_211 <= c_reg_210 | data_from_out_mat_13_3;
      c_reg_212 <= c_reg_211 | data_from_out_mat_13_4;
      c_reg_213 <= c_reg_212 | data_from_out_mat_13_5;
      c_reg_214 <= c_reg_213 | data_from_out_mat_13_6;
      c_reg_215 <= c_reg_214 | data_from_out_mat_13_7;
      c_reg_216 <= c_reg_215 | data_from_out_mat_13_8;
      c_reg_217 <= c_reg_216 | data_from_out_mat_13_9;
      c_reg_218 <= c_reg_217 | data_from_out_mat_13_10;
      c_reg_219 <= c_reg_218 | data_from_out_mat_13_11;
      c_reg_220 <= c_reg_219 | data_from_out_mat_13_12;
      c_reg_221 <= c_reg_220 | data_from_out_mat_13_13;
      c_reg_222 <= c_reg_221 | data_from_out_mat_13_14;
      c_reg_223 <= c_reg_222 | data_from_out_mat_13_15;
      c_reg_224 <= c_reg_223 | data_from_out_mat_14_0;
      c_reg_225 <= c_reg_224 | data_from_out_mat_14_1;
      c_reg_226 <= c_reg_225 | data_from_out_mat_14_2;
      c_reg_227 <= c_reg_226 | data_from_out_mat_14_3;
      c_reg_228 <= c_reg_227 | data_from_out_mat_14_4;
      c_reg_229 <= c_reg_228 | data_from_out_mat_14_5;
      c_reg_230 <= c_reg_229 | data_from_out_mat_14_6;
      c_reg_231 <= c_reg_230 | data_from_out_mat_14_7;
      c_reg_232 <= c_reg_231 | data_from_out_mat_14_8;
      c_reg_233 <= c_reg_232 | data_from_out_mat_14_9;
      c_reg_234 <= c_reg_233 | data_from_out_mat_14_10;
      c_reg_235 <= c_reg_234 | data_from_out_mat_14_11;
      c_reg_236 <= c_reg_235 | data_from_out_mat_14_12;
      c_reg_237 <= c_reg_236 | data_from_out_mat_14_13;
      c_reg_238 <= c_reg_237 | data_from_out_mat_14_14;
      c_reg_239 <= c_reg_238 | data_from_out_mat_14_15;
      c_reg_240 <= c_reg_239 | data_from_out_mat_15_0;
      c_reg_241 <= c_reg_240 | data_from_out_mat_15_1;
      c_reg_242 <= c_reg_241 | data_from_out_mat_15_2;
      c_reg_243 <= c_reg_242 | data_from_out_mat_15_3;
      c_reg_244 <= c_reg_243 | data_from_out_mat_15_4;
      c_reg_245 <= c_reg_244 | data_from_out_mat_15_5;
      c_reg_246 <= c_reg_245 | data_from_out_mat_15_6;
      c_reg_247 <= c_reg_246 | data_from_out_mat_15_7;
      c_reg_248 <= c_reg_247 | data_from_out_mat_15_8;
      c_reg_249 <= c_reg_248 | data_from_out_mat_15_9;
      c_reg_250 <= c_reg_249 | data_from_out_mat_15_10;
      c_reg_251 <= c_reg_250 | data_from_out_mat_15_11;
      c_reg_252 <= c_reg_251 | data_from_out_mat_15_12;
      c_reg_253 <= c_reg_252 | data_from_out_mat_15_13;
      c_reg_254 <= c_reg_253 | data_from_out_mat_15_14;
      c_reg_255 <= c_reg_254 | data_from_out_mat_15_15;
      data_from_out_mat <= c_reg_255;
    end
  end

  //  BRAM matrix C0_0
  ram matrix_c_0_0 (
    .addr0(c_addr_muxed_0_0_reg),
    .d0(c_data_0_0),
    .we0(we_c),
    .q0(data_from_out_mat_0_0),
    .clk(clk));

  //  BRAM matrix C0_1
  ram matrix_c_0_1 (
    .addr0(c_addr_muxed_0_1_reg),
    .d0(c_data_0_1),
    .we0(we_c),
    .q0(data_from_out_mat_0_1),
    .clk(clk));

  //  BRAM matrix C0_2
  ram matrix_c_0_2 (
    .addr0(c_addr_muxed_0_2_reg),
    .d0(c_data_0_2),
    .we0(we_c),
    .q0(data_from_out_mat_0_2),
    .clk(clk));

  //  BRAM matrix C0_3
  ram matrix_c_0_3 (
    .addr0(c_addr_muxed_0_3_reg),
    .d0(c_data_0_3),
    .we0(we_c),
    .q0(data_from_out_mat_0_3),
    .clk(clk));

  //  BRAM matrix C0_4
  ram matrix_c_0_4 (
    .addr0(c_addr_muxed_0_4_reg),
    .d0(c_data_0_4),
    .we0(we_c),
    .q0(data_from_out_mat_0_4),
    .clk(clk));

  //  BRAM matrix C0_5
  ram matrix_c_0_5 (
    .addr0(c_addr_muxed_0_5_reg),
    .d0(c_data_0_5),
    .we0(we_c),
    .q0(data_from_out_mat_0_5),
    .clk(clk));

  //  BRAM matrix C0_6
  ram matrix_c_0_6 (
    .addr0(c_addr_muxed_0_6_reg),
    .d0(c_data_0_6),
    .we0(we_c),
    .q0(data_from_out_mat_0_6),
    .clk(clk));

  //  BRAM matrix C0_7
  ram matrix_c_0_7 (
    .addr0(c_addr_muxed_0_7_reg),
    .d0(c_data_0_7),
    .we0(we_c),
    .q0(data_from_out_mat_0_7),
    .clk(clk));

  //  BRAM matrix C0_8
  ram matrix_c_0_8 (
    .addr0(c_addr_muxed_0_8_reg),
    .d0(c_data_0_8),
    .we0(we_c),
    .q0(data_from_out_mat_0_8),
    .clk(clk));

  //  BRAM matrix C0_9
  ram matrix_c_0_9 (
    .addr0(c_addr_muxed_0_9_reg),
    .d0(c_data_0_9),
    .we0(we_c),
    .q0(data_from_out_mat_0_9),
    .clk(clk));

  //  BRAM matrix C0_10
  ram matrix_c_0_10 (
    .addr0(c_addr_muxed_0_10_reg),
    .d0(c_data_0_10),
    .we0(we_c),
    .q0(data_from_out_mat_0_10),
    .clk(clk));

  //  BRAM matrix C0_11
  ram matrix_c_0_11 (
    .addr0(c_addr_muxed_0_11_reg),
    .d0(c_data_0_11),
    .we0(we_c),
    .q0(data_from_out_mat_0_11),
    .clk(clk));

  //  BRAM matrix C0_12
  ram matrix_c_0_12 (
    .addr0(c_addr_muxed_0_12_reg),
    .d0(c_data_0_12),
    .we0(we_c),
    .q0(data_from_out_mat_0_12),
    .clk(clk));

  //  BRAM matrix C0_13
  ram matrix_c_0_13 (
    .addr0(c_addr_muxed_0_13_reg),
    .d0(c_data_0_13),
    .we0(we_c),
    .q0(data_from_out_mat_0_13),
    .clk(clk));

  //  BRAM matrix C0_14
  ram matrix_c_0_14 (
    .addr0(c_addr_muxed_0_14_reg),
    .d0(c_data_0_14),
    .we0(we_c),
    .q0(data_from_out_mat_0_14),
    .clk(clk));

  //  BRAM matrix C0_15
  ram matrix_c_0_15 (
    .addr0(c_addr_muxed_0_15_reg),
    .d0(c_data_0_15),
    .we0(we_c),
    .q0(data_from_out_mat_0_15),
    .clk(clk));

  //  BRAM matrix C1_0
  ram matrix_c_1_0 (
    .addr0(c_addr_muxed_1_0_reg),
    .d0(c_data_1_0),
    .we0(we_c),
    .q0(data_from_out_mat_1_0),
    .clk(clk));

  //  BRAM matrix C1_1
  ram matrix_c_1_1 (
    .addr0(c_addr_muxed_1_1_reg),
    .d0(c_data_1_1),
    .we0(we_c),
    .q0(data_from_out_mat_1_1),
    .clk(clk));

  //  BRAM matrix C1_2
  ram matrix_c_1_2 (
    .addr0(c_addr_muxed_1_2_reg),
    .d0(c_data_1_2),
    .we0(we_c),
    .q0(data_from_out_mat_1_2),
    .clk(clk));

  //  BRAM matrix C1_3
  ram matrix_c_1_3 (
    .addr0(c_addr_muxed_1_3_reg),
    .d0(c_data_1_3),
    .we0(we_c),
    .q0(data_from_out_mat_1_3),
    .clk(clk));

  //  BRAM matrix C1_4
  ram matrix_c_1_4 (
    .addr0(c_addr_muxed_1_4_reg),
    .d0(c_data_1_4),
    .we0(we_c),
    .q0(data_from_out_mat_1_4),
    .clk(clk));

  //  BRAM matrix C1_5
  ram matrix_c_1_5 (
    .addr0(c_addr_muxed_1_5_reg),
    .d0(c_data_1_5),
    .we0(we_c),
    .q0(data_from_out_mat_1_5),
    .clk(clk));

  //  BRAM matrix C1_6
  ram matrix_c_1_6 (
    .addr0(c_addr_muxed_1_6_reg),
    .d0(c_data_1_6),
    .we0(we_c),
    .q0(data_from_out_mat_1_6),
    .clk(clk));

  //  BRAM matrix C1_7
  ram matrix_c_1_7 (
    .addr0(c_addr_muxed_1_7_reg),
    .d0(c_data_1_7),
    .we0(we_c),
    .q0(data_from_out_mat_1_7),
    .clk(clk));

  //  BRAM matrix C1_8
  ram matrix_c_1_8 (
    .addr0(c_addr_muxed_1_8_reg),
    .d0(c_data_1_8),
    .we0(we_c),
    .q0(data_from_out_mat_1_8),
    .clk(clk));

  //  BRAM matrix C1_9
  ram matrix_c_1_9 (
    .addr0(c_addr_muxed_1_9_reg),
    .d0(c_data_1_9),
    .we0(we_c),
    .q0(data_from_out_mat_1_9),
    .clk(clk));

  //  BRAM matrix C1_10
  ram matrix_c_1_10 (
    .addr0(c_addr_muxed_1_10_reg),
    .d0(c_data_1_10),
    .we0(we_c),
    .q0(data_from_out_mat_1_10),
    .clk(clk));

  //  BRAM matrix C1_11
  ram matrix_c_1_11 (
    .addr0(c_addr_muxed_1_11_reg),
    .d0(c_data_1_11),
    .we0(we_c),
    .q0(data_from_out_mat_1_11),
    .clk(clk));

  //  BRAM matrix C1_12
  ram matrix_c_1_12 (
    .addr0(c_addr_muxed_1_12_reg),
    .d0(c_data_1_12),
    .we0(we_c),
    .q0(data_from_out_mat_1_12),
    .clk(clk));

  //  BRAM matrix C1_13
  ram matrix_c_1_13 (
    .addr0(c_addr_muxed_1_13_reg),
    .d0(c_data_1_13),
    .we0(we_c),
    .q0(data_from_out_mat_1_13),
    .clk(clk));

  //  BRAM matrix C1_14
  ram matrix_c_1_14 (
    .addr0(c_addr_muxed_1_14_reg),
    .d0(c_data_1_14),
    .we0(we_c),
    .q0(data_from_out_mat_1_14),
    .clk(clk));

  //  BRAM matrix C1_15
  ram matrix_c_1_15 (
    .addr0(c_addr_muxed_1_15_reg),
    .d0(c_data_1_15),
    .we0(we_c),
    .q0(data_from_out_mat_1_15),
    .clk(clk));

  //  BRAM matrix C2_0
  ram matrix_c_2_0 (
    .addr0(c_addr_muxed_2_0_reg),
    .d0(c_data_2_0),
    .we0(we_c),
    .q0(data_from_out_mat_2_0),
    .clk(clk));

  //  BRAM matrix C2_1
  ram matrix_c_2_1 (
    .addr0(c_addr_muxed_2_1_reg),
    .d0(c_data_2_1),
    .we0(we_c),
    .q0(data_from_out_mat_2_1),
    .clk(clk));

  //  BRAM matrix C2_2
  ram matrix_c_2_2 (
    .addr0(c_addr_muxed_2_2_reg),
    .d0(c_data_2_2),
    .we0(we_c),
    .q0(data_from_out_mat_2_2),
    .clk(clk));

  //  BRAM matrix C2_3
  ram matrix_c_2_3 (
    .addr0(c_addr_muxed_2_3_reg),
    .d0(c_data_2_3),
    .we0(we_c),
    .q0(data_from_out_mat_2_3),
    .clk(clk));

  //  BRAM matrix C2_4
  ram matrix_c_2_4 (
    .addr0(c_addr_muxed_2_4_reg),
    .d0(c_data_2_4),
    .we0(we_c),
    .q0(data_from_out_mat_2_4),
    .clk(clk));

  //  BRAM matrix C2_5
  ram matrix_c_2_5 (
    .addr0(c_addr_muxed_2_5_reg),
    .d0(c_data_2_5),
    .we0(we_c),
    .q0(data_from_out_mat_2_5),
    .clk(clk));

  //  BRAM matrix C2_6
  ram matrix_c_2_6 (
    .addr0(c_addr_muxed_2_6_reg),
    .d0(c_data_2_6),
    .we0(we_c),
    .q0(data_from_out_mat_2_6),
    .clk(clk));

  //  BRAM matrix C2_7
  ram matrix_c_2_7 (
    .addr0(c_addr_muxed_2_7_reg),
    .d0(c_data_2_7),
    .we0(we_c),
    .q0(data_from_out_mat_2_7),
    .clk(clk));

  //  BRAM matrix C2_8
  ram matrix_c_2_8 (
    .addr0(c_addr_muxed_2_8_reg),
    .d0(c_data_2_8),
    .we0(we_c),
    .q0(data_from_out_mat_2_8),
    .clk(clk));

  //  BRAM matrix C2_9
  ram matrix_c_2_9 (
    .addr0(c_addr_muxed_2_9_reg),
    .d0(c_data_2_9),
    .we0(we_c),
    .q0(data_from_out_mat_2_9),
    .clk(clk));

  //  BRAM matrix C2_10
  ram matrix_c_2_10 (
    .addr0(c_addr_muxed_2_10_reg),
    .d0(c_data_2_10),
    .we0(we_c),
    .q0(data_from_out_mat_2_10),
    .clk(clk));

  //  BRAM matrix C2_11
  ram matrix_c_2_11 (
    .addr0(c_addr_muxed_2_11_reg),
    .d0(c_data_2_11),
    .we0(we_c),
    .q0(data_from_out_mat_2_11),
    .clk(clk));

  //  BRAM matrix C2_12
  ram matrix_c_2_12 (
    .addr0(c_addr_muxed_2_12_reg),
    .d0(c_data_2_12),
    .we0(we_c),
    .q0(data_from_out_mat_2_12),
    .clk(clk));

  //  BRAM matrix C2_13
  ram matrix_c_2_13 (
    .addr0(c_addr_muxed_2_13_reg),
    .d0(c_data_2_13),
    .we0(we_c),
    .q0(data_from_out_mat_2_13),
    .clk(clk));

  //  BRAM matrix C2_14
  ram matrix_c_2_14 (
    .addr0(c_addr_muxed_2_14_reg),
    .d0(c_data_2_14),
    .we0(we_c),
    .q0(data_from_out_mat_2_14),
    .clk(clk));

  //  BRAM matrix C2_15
  ram matrix_c_2_15 (
    .addr0(c_addr_muxed_2_15_reg),
    .d0(c_data_2_15),
    .we0(we_c),
    .q0(data_from_out_mat_2_15),
    .clk(clk));

  //  BRAM matrix C3_0
  ram matrix_c_3_0 (
    .addr0(c_addr_muxed_3_0_reg),
    .d0(c_data_3_0),
    .we0(we_c),
    .q0(data_from_out_mat_3_0),
    .clk(clk));

  //  BRAM matrix C3_1
  ram matrix_c_3_1 (
    .addr0(c_addr_muxed_3_1_reg),
    .d0(c_data_3_1),
    .we0(we_c),
    .q0(data_from_out_mat_3_1),
    .clk(clk));

  //  BRAM matrix C3_2
  ram matrix_c_3_2 (
    .addr0(c_addr_muxed_3_2_reg),
    .d0(c_data_3_2),
    .we0(we_c),
    .q0(data_from_out_mat_3_2),
    .clk(clk));

  //  BRAM matrix C3_3
  ram matrix_c_3_3 (
    .addr0(c_addr_muxed_3_3_reg),
    .d0(c_data_3_3),
    .we0(we_c),
    .q0(data_from_out_mat_3_3),
    .clk(clk));

  //  BRAM matrix C3_4
  ram matrix_c_3_4 (
    .addr0(c_addr_muxed_3_4_reg),
    .d0(c_data_3_4),
    .we0(we_c),
    .q0(data_from_out_mat_3_4),
    .clk(clk));

  //  BRAM matrix C3_5
  ram matrix_c_3_5 (
    .addr0(c_addr_muxed_3_5_reg),
    .d0(c_data_3_5),
    .we0(we_c),
    .q0(data_from_out_mat_3_5),
    .clk(clk));

  //  BRAM matrix C3_6
  ram matrix_c_3_6 (
    .addr0(c_addr_muxed_3_6_reg),
    .d0(c_data_3_6),
    .we0(we_c),
    .q0(data_from_out_mat_3_6),
    .clk(clk));

  //  BRAM matrix C3_7
  ram matrix_c_3_7 (
    .addr0(c_addr_muxed_3_7_reg),
    .d0(c_data_3_7),
    .we0(we_c),
    .q0(data_from_out_mat_3_7),
    .clk(clk));

  //  BRAM matrix C3_8
  ram matrix_c_3_8 (
    .addr0(c_addr_muxed_3_8_reg),
    .d0(c_data_3_8),
    .we0(we_c),
    .q0(data_from_out_mat_3_8),
    .clk(clk));

  //  BRAM matrix C3_9
  ram matrix_c_3_9 (
    .addr0(c_addr_muxed_3_9_reg),
    .d0(c_data_3_9),
    .we0(we_c),
    .q0(data_from_out_mat_3_9),
    .clk(clk));

  //  BRAM matrix C3_10
  ram matrix_c_3_10 (
    .addr0(c_addr_muxed_3_10_reg),
    .d0(c_data_3_10),
    .we0(we_c),
    .q0(data_from_out_mat_3_10),
    .clk(clk));

  //  BRAM matrix C3_11
  ram matrix_c_3_11 (
    .addr0(c_addr_muxed_3_11_reg),
    .d0(c_data_3_11),
    .we0(we_c),
    .q0(data_from_out_mat_3_11),
    .clk(clk));

  //  BRAM matrix C3_12
  ram matrix_c_3_12 (
    .addr0(c_addr_muxed_3_12_reg),
    .d0(c_data_3_12),
    .we0(we_c),
    .q0(data_from_out_mat_3_12),
    .clk(clk));

  //  BRAM matrix C3_13
  ram matrix_c_3_13 (
    .addr0(c_addr_muxed_3_13_reg),
    .d0(c_data_3_13),
    .we0(we_c),
    .q0(data_from_out_mat_3_13),
    .clk(clk));

  //  BRAM matrix C3_14
  ram matrix_c_3_14 (
    .addr0(c_addr_muxed_3_14_reg),
    .d0(c_data_3_14),
    .we0(we_c),
    .q0(data_from_out_mat_3_14),
    .clk(clk));

  //  BRAM matrix C3_15
  ram matrix_c_3_15 (
    .addr0(c_addr_muxed_3_15_reg),
    .d0(c_data_3_15),
    .we0(we_c),
    .q0(data_from_out_mat_3_15),
    .clk(clk));

  //  BRAM matrix C4_0
  ram matrix_c_4_0 (
    .addr0(c_addr_muxed_4_0_reg),
    .d0(c_data_4_0),
    .we0(we_c),
    .q0(data_from_out_mat_4_0),
    .clk(clk));

  //  BRAM matrix C4_1
  ram matrix_c_4_1 (
    .addr0(c_addr_muxed_4_1_reg),
    .d0(c_data_4_1),
    .we0(we_c),
    .q0(data_from_out_mat_4_1),
    .clk(clk));

  //  BRAM matrix C4_2
  ram matrix_c_4_2 (
    .addr0(c_addr_muxed_4_2_reg),
    .d0(c_data_4_2),
    .we0(we_c),
    .q0(data_from_out_mat_4_2),
    .clk(clk));

  //  BRAM matrix C4_3
  ram matrix_c_4_3 (
    .addr0(c_addr_muxed_4_3_reg),
    .d0(c_data_4_3),
    .we0(we_c),
    .q0(data_from_out_mat_4_3),
    .clk(clk));

  //  BRAM matrix C4_4
  ram matrix_c_4_4 (
    .addr0(c_addr_muxed_4_4_reg),
    .d0(c_data_4_4),
    .we0(we_c),
    .q0(data_from_out_mat_4_4),
    .clk(clk));

  //  BRAM matrix C4_5
  ram matrix_c_4_5 (
    .addr0(c_addr_muxed_4_5_reg),
    .d0(c_data_4_5),
    .we0(we_c),
    .q0(data_from_out_mat_4_5),
    .clk(clk));

  //  BRAM matrix C4_6
  ram matrix_c_4_6 (
    .addr0(c_addr_muxed_4_6_reg),
    .d0(c_data_4_6),
    .we0(we_c),
    .q0(data_from_out_mat_4_6),
    .clk(clk));

  //  BRAM matrix C4_7
  ram matrix_c_4_7 (
    .addr0(c_addr_muxed_4_7_reg),
    .d0(c_data_4_7),
    .we0(we_c),
    .q0(data_from_out_mat_4_7),
    .clk(clk));

  //  BRAM matrix C4_8
  ram matrix_c_4_8 (
    .addr0(c_addr_muxed_4_8_reg),
    .d0(c_data_4_8),
    .we0(we_c),
    .q0(data_from_out_mat_4_8),
    .clk(clk));

  //  BRAM matrix C4_9
  ram matrix_c_4_9 (
    .addr0(c_addr_muxed_4_9_reg),
    .d0(c_data_4_9),
    .we0(we_c),
    .q0(data_from_out_mat_4_9),
    .clk(clk));

  //  BRAM matrix C4_10
  ram matrix_c_4_10 (
    .addr0(c_addr_muxed_4_10_reg),
    .d0(c_data_4_10),
    .we0(we_c),
    .q0(data_from_out_mat_4_10),
    .clk(clk));

  //  BRAM matrix C4_11
  ram matrix_c_4_11 (
    .addr0(c_addr_muxed_4_11_reg),
    .d0(c_data_4_11),
    .we0(we_c),
    .q0(data_from_out_mat_4_11),
    .clk(clk));

  //  BRAM matrix C4_12
  ram matrix_c_4_12 (
    .addr0(c_addr_muxed_4_12_reg),
    .d0(c_data_4_12),
    .we0(we_c),
    .q0(data_from_out_mat_4_12),
    .clk(clk));

  //  BRAM matrix C4_13
  ram matrix_c_4_13 (
    .addr0(c_addr_muxed_4_13_reg),
    .d0(c_data_4_13),
    .we0(we_c),
    .q0(data_from_out_mat_4_13),
    .clk(clk));

  //  BRAM matrix C4_14
  ram matrix_c_4_14 (
    .addr0(c_addr_muxed_4_14_reg),
    .d0(c_data_4_14),
    .we0(we_c),
    .q0(data_from_out_mat_4_14),
    .clk(clk));

  //  BRAM matrix C4_15
  ram matrix_c_4_15 (
    .addr0(c_addr_muxed_4_15_reg),
    .d0(c_data_4_15),
    .we0(we_c),
    .q0(data_from_out_mat_4_15),
    .clk(clk));

  //  BRAM matrix C5_0
  ram matrix_c_5_0 (
    .addr0(c_addr_muxed_5_0_reg),
    .d0(c_data_5_0),
    .we0(we_c),
    .q0(data_from_out_mat_5_0),
    .clk(clk));

  //  BRAM matrix C5_1
  ram matrix_c_5_1 (
    .addr0(c_addr_muxed_5_1_reg),
    .d0(c_data_5_1),
    .we0(we_c),
    .q0(data_from_out_mat_5_1),
    .clk(clk));

  //  BRAM matrix C5_2
  ram matrix_c_5_2 (
    .addr0(c_addr_muxed_5_2_reg),
    .d0(c_data_5_2),
    .we0(we_c),
    .q0(data_from_out_mat_5_2),
    .clk(clk));

  //  BRAM matrix C5_3
  ram matrix_c_5_3 (
    .addr0(c_addr_muxed_5_3_reg),
    .d0(c_data_5_3),
    .we0(we_c),
    .q0(data_from_out_mat_5_3),
    .clk(clk));

  //  BRAM matrix C5_4
  ram matrix_c_5_4 (
    .addr0(c_addr_muxed_5_4_reg),
    .d0(c_data_5_4),
    .we0(we_c),
    .q0(data_from_out_mat_5_4),
    .clk(clk));

  //  BRAM matrix C5_5
  ram matrix_c_5_5 (
    .addr0(c_addr_muxed_5_5_reg),
    .d0(c_data_5_5),
    .we0(we_c),
    .q0(data_from_out_mat_5_5),
    .clk(clk));

  //  BRAM matrix C5_6
  ram matrix_c_5_6 (
    .addr0(c_addr_muxed_5_6_reg),
    .d0(c_data_5_6),
    .we0(we_c),
    .q0(data_from_out_mat_5_6),
    .clk(clk));

  //  BRAM matrix C5_7
  ram matrix_c_5_7 (
    .addr0(c_addr_muxed_5_7_reg),
    .d0(c_data_5_7),
    .we0(we_c),
    .q0(data_from_out_mat_5_7),
    .clk(clk));

  //  BRAM matrix C5_8
  ram matrix_c_5_8 (
    .addr0(c_addr_muxed_5_8_reg),
    .d0(c_data_5_8),
    .we0(we_c),
    .q0(data_from_out_mat_5_8),
    .clk(clk));

  //  BRAM matrix C5_9
  ram matrix_c_5_9 (
    .addr0(c_addr_muxed_5_9_reg),
    .d0(c_data_5_9),
    .we0(we_c),
    .q0(data_from_out_mat_5_9),
    .clk(clk));

  //  BRAM matrix C5_10
  ram matrix_c_5_10 (
    .addr0(c_addr_muxed_5_10_reg),
    .d0(c_data_5_10),
    .we0(we_c),
    .q0(data_from_out_mat_5_10),
    .clk(clk));

  //  BRAM matrix C5_11
  ram matrix_c_5_11 (
    .addr0(c_addr_muxed_5_11_reg),
    .d0(c_data_5_11),
    .we0(we_c),
    .q0(data_from_out_mat_5_11),
    .clk(clk));

  //  BRAM matrix C5_12
  ram matrix_c_5_12 (
    .addr0(c_addr_muxed_5_12_reg),
    .d0(c_data_5_12),
    .we0(we_c),
    .q0(data_from_out_mat_5_12),
    .clk(clk));

  //  BRAM matrix C5_13
  ram matrix_c_5_13 (
    .addr0(c_addr_muxed_5_13_reg),
    .d0(c_data_5_13),
    .we0(we_c),
    .q0(data_from_out_mat_5_13),
    .clk(clk));

  //  BRAM matrix C5_14
  ram matrix_c_5_14 (
    .addr0(c_addr_muxed_5_14_reg),
    .d0(c_data_5_14),
    .we0(we_c),
    .q0(data_from_out_mat_5_14),
    .clk(clk));

  //  BRAM matrix C5_15
  ram matrix_c_5_15 (
    .addr0(c_addr_muxed_5_15_reg),
    .d0(c_data_5_15),
    .we0(we_c),
    .q0(data_from_out_mat_5_15),
    .clk(clk));

  //  BRAM matrix C6_0
  ram matrix_c_6_0 (
    .addr0(c_addr_muxed_6_0_reg),
    .d0(c_data_6_0),
    .we0(we_c),
    .q0(data_from_out_mat_6_0),
    .clk(clk));

  //  BRAM matrix C6_1
  ram matrix_c_6_1 (
    .addr0(c_addr_muxed_6_1_reg),
    .d0(c_data_6_1),
    .we0(we_c),
    .q0(data_from_out_mat_6_1),
    .clk(clk));

  //  BRAM matrix C6_2
  ram matrix_c_6_2 (
    .addr0(c_addr_muxed_6_2_reg),
    .d0(c_data_6_2),
    .we0(we_c),
    .q0(data_from_out_mat_6_2),
    .clk(clk));

  //  BRAM matrix C6_3
  ram matrix_c_6_3 (
    .addr0(c_addr_muxed_6_3_reg),
    .d0(c_data_6_3),
    .we0(we_c),
    .q0(data_from_out_mat_6_3),
    .clk(clk));

  //  BRAM matrix C6_4
  ram matrix_c_6_4 (
    .addr0(c_addr_muxed_6_4_reg),
    .d0(c_data_6_4),
    .we0(we_c),
    .q0(data_from_out_mat_6_4),
    .clk(clk));

  //  BRAM matrix C6_5
  ram matrix_c_6_5 (
    .addr0(c_addr_muxed_6_5_reg),
    .d0(c_data_6_5),
    .we0(we_c),
    .q0(data_from_out_mat_6_5),
    .clk(clk));

  //  BRAM matrix C6_6
  ram matrix_c_6_6 (
    .addr0(c_addr_muxed_6_6_reg),
    .d0(c_data_6_6),
    .we0(we_c),
    .q0(data_from_out_mat_6_6),
    .clk(clk));

  //  BRAM matrix C6_7
  ram matrix_c_6_7 (
    .addr0(c_addr_muxed_6_7_reg),
    .d0(c_data_6_7),
    .we0(we_c),
    .q0(data_from_out_mat_6_7),
    .clk(clk));

  //  BRAM matrix C6_8
  ram matrix_c_6_8 (
    .addr0(c_addr_muxed_6_8_reg),
    .d0(c_data_6_8),
    .we0(we_c),
    .q0(data_from_out_mat_6_8),
    .clk(clk));

  //  BRAM matrix C6_9
  ram matrix_c_6_9 (
    .addr0(c_addr_muxed_6_9_reg),
    .d0(c_data_6_9),
    .we0(we_c),
    .q0(data_from_out_mat_6_9),
    .clk(clk));

  //  BRAM matrix C6_10
  ram matrix_c_6_10 (
    .addr0(c_addr_muxed_6_10_reg),
    .d0(c_data_6_10),
    .we0(we_c),
    .q0(data_from_out_mat_6_10),
    .clk(clk));

  //  BRAM matrix C6_11
  ram matrix_c_6_11 (
    .addr0(c_addr_muxed_6_11_reg),
    .d0(c_data_6_11),
    .we0(we_c),
    .q0(data_from_out_mat_6_11),
    .clk(clk));

  //  BRAM matrix C6_12
  ram matrix_c_6_12 (
    .addr0(c_addr_muxed_6_12_reg),
    .d0(c_data_6_12),
    .we0(we_c),
    .q0(data_from_out_mat_6_12),
    .clk(clk));

  //  BRAM matrix C6_13
  ram matrix_c_6_13 (
    .addr0(c_addr_muxed_6_13_reg),
    .d0(c_data_6_13),
    .we0(we_c),
    .q0(data_from_out_mat_6_13),
    .clk(clk));

  //  BRAM matrix C6_14
  ram matrix_c_6_14 (
    .addr0(c_addr_muxed_6_14_reg),
    .d0(c_data_6_14),
    .we0(we_c),
    .q0(data_from_out_mat_6_14),
    .clk(clk));

  //  BRAM matrix C6_15
  ram matrix_c_6_15 (
    .addr0(c_addr_muxed_6_15_reg),
    .d0(c_data_6_15),
    .we0(we_c),
    .q0(data_from_out_mat_6_15),
    .clk(clk));

  //  BRAM matrix C7_0
  ram matrix_c_7_0 (
    .addr0(c_addr_muxed_7_0_reg),
    .d0(c_data_7_0),
    .we0(we_c),
    .q0(data_from_out_mat_7_0),
    .clk(clk));

  //  BRAM matrix C7_1
  ram matrix_c_7_1 (
    .addr0(c_addr_muxed_7_1_reg),
    .d0(c_data_7_1),
    .we0(we_c),
    .q0(data_from_out_mat_7_1),
    .clk(clk));

  //  BRAM matrix C7_2
  ram matrix_c_7_2 (
    .addr0(c_addr_muxed_7_2_reg),
    .d0(c_data_7_2),
    .we0(we_c),
    .q0(data_from_out_mat_7_2),
    .clk(clk));

  //  BRAM matrix C7_3
  ram matrix_c_7_3 (
    .addr0(c_addr_muxed_7_3_reg),
    .d0(c_data_7_3),
    .we0(we_c),
    .q0(data_from_out_mat_7_3),
    .clk(clk));

  //  BRAM matrix C7_4
  ram matrix_c_7_4 (
    .addr0(c_addr_muxed_7_4_reg),
    .d0(c_data_7_4),
    .we0(we_c),
    .q0(data_from_out_mat_7_4),
    .clk(clk));

  //  BRAM matrix C7_5
  ram matrix_c_7_5 (
    .addr0(c_addr_muxed_7_5_reg),
    .d0(c_data_7_5),
    .we0(we_c),
    .q0(data_from_out_mat_7_5),
    .clk(clk));

  //  BRAM matrix C7_6
  ram matrix_c_7_6 (
    .addr0(c_addr_muxed_7_6_reg),
    .d0(c_data_7_6),
    .we0(we_c),
    .q0(data_from_out_mat_7_6),
    .clk(clk));

  //  BRAM matrix C7_7
  ram matrix_c_7_7 (
    .addr0(c_addr_muxed_7_7_reg),
    .d0(c_data_7_7),
    .we0(we_c),
    .q0(data_from_out_mat_7_7),
    .clk(clk));

  //  BRAM matrix C7_8
  ram matrix_c_7_8 (
    .addr0(c_addr_muxed_7_8_reg),
    .d0(c_data_7_8),
    .we0(we_c),
    .q0(data_from_out_mat_7_8),
    .clk(clk));

  //  BRAM matrix C7_9
  ram matrix_c_7_9 (
    .addr0(c_addr_muxed_7_9_reg),
    .d0(c_data_7_9),
    .we0(we_c),
    .q0(data_from_out_mat_7_9),
    .clk(clk));

  //  BRAM matrix C7_10
  ram matrix_c_7_10 (
    .addr0(c_addr_muxed_7_10_reg),
    .d0(c_data_7_10),
    .we0(we_c),
    .q0(data_from_out_mat_7_10),
    .clk(clk));

  //  BRAM matrix C7_11
  ram matrix_c_7_11 (
    .addr0(c_addr_muxed_7_11_reg),
    .d0(c_data_7_11),
    .we0(we_c),
    .q0(data_from_out_mat_7_11),
    .clk(clk));

  //  BRAM matrix C7_12
  ram matrix_c_7_12 (
    .addr0(c_addr_muxed_7_12_reg),
    .d0(c_data_7_12),
    .we0(we_c),
    .q0(data_from_out_mat_7_12),
    .clk(clk));

  //  BRAM matrix C7_13
  ram matrix_c_7_13 (
    .addr0(c_addr_muxed_7_13_reg),
    .d0(c_data_7_13),
    .we0(we_c),
    .q0(data_from_out_mat_7_13),
    .clk(clk));

  //  BRAM matrix C7_14
  ram matrix_c_7_14 (
    .addr0(c_addr_muxed_7_14_reg),
    .d0(c_data_7_14),
    .we0(we_c),
    .q0(data_from_out_mat_7_14),
    .clk(clk));

  //  BRAM matrix C7_15
  ram matrix_c_7_15 (
    .addr0(c_addr_muxed_7_15_reg),
    .d0(c_data_7_15),
    .we0(we_c),
    .q0(data_from_out_mat_7_15),
    .clk(clk));

  //  BRAM matrix C8_0
  ram matrix_c_8_0 (
    .addr0(c_addr_muxed_8_0_reg),
    .d0(c_data_8_0),
    .we0(we_c),
    .q0(data_from_out_mat_8_0),
    .clk(clk));

  //  BRAM matrix C8_1
  ram matrix_c_8_1 (
    .addr0(c_addr_muxed_8_1_reg),
    .d0(c_data_8_1),
    .we0(we_c),
    .q0(data_from_out_mat_8_1),
    .clk(clk));

  //  BRAM matrix C8_2
  ram matrix_c_8_2 (
    .addr0(c_addr_muxed_8_2_reg),
    .d0(c_data_8_2),
    .we0(we_c),
    .q0(data_from_out_mat_8_2),
    .clk(clk));

  //  BRAM matrix C8_3
  ram matrix_c_8_3 (
    .addr0(c_addr_muxed_8_3_reg),
    .d0(c_data_8_3),
    .we0(we_c),
    .q0(data_from_out_mat_8_3),
    .clk(clk));

  //  BRAM matrix C8_4
  ram matrix_c_8_4 (
    .addr0(c_addr_muxed_8_4_reg),
    .d0(c_data_8_4),
    .we0(we_c),
    .q0(data_from_out_mat_8_4),
    .clk(clk));

  //  BRAM matrix C8_5
  ram matrix_c_8_5 (
    .addr0(c_addr_muxed_8_5_reg),
    .d0(c_data_8_5),
    .we0(we_c),
    .q0(data_from_out_mat_8_5),
    .clk(clk));

  //  BRAM matrix C8_6
  ram matrix_c_8_6 (
    .addr0(c_addr_muxed_8_6_reg),
    .d0(c_data_8_6),
    .we0(we_c),
    .q0(data_from_out_mat_8_6),
    .clk(clk));

  //  BRAM matrix C8_7
  ram matrix_c_8_7 (
    .addr0(c_addr_muxed_8_7_reg),
    .d0(c_data_8_7),
    .we0(we_c),
    .q0(data_from_out_mat_8_7),
    .clk(clk));

  //  BRAM matrix C8_8
  ram matrix_c_8_8 (
    .addr0(c_addr_muxed_8_8_reg),
    .d0(c_data_8_8),
    .we0(we_c),
    .q0(data_from_out_mat_8_8),
    .clk(clk));

  //  BRAM matrix C8_9
  ram matrix_c_8_9 (
    .addr0(c_addr_muxed_8_9_reg),
    .d0(c_data_8_9),
    .we0(we_c),
    .q0(data_from_out_mat_8_9),
    .clk(clk));

  //  BRAM matrix C8_10
  ram matrix_c_8_10 (
    .addr0(c_addr_muxed_8_10_reg),
    .d0(c_data_8_10),
    .we0(we_c),
    .q0(data_from_out_mat_8_10),
    .clk(clk));

  //  BRAM matrix C8_11
  ram matrix_c_8_11 (
    .addr0(c_addr_muxed_8_11_reg),
    .d0(c_data_8_11),
    .we0(we_c),
    .q0(data_from_out_mat_8_11),
    .clk(clk));

  //  BRAM matrix C8_12
  ram matrix_c_8_12 (
    .addr0(c_addr_muxed_8_12_reg),
    .d0(c_data_8_12),
    .we0(we_c),
    .q0(data_from_out_mat_8_12),
    .clk(clk));

  //  BRAM matrix C8_13
  ram matrix_c_8_13 (
    .addr0(c_addr_muxed_8_13_reg),
    .d0(c_data_8_13),
    .we0(we_c),
    .q0(data_from_out_mat_8_13),
    .clk(clk));

  //  BRAM matrix C8_14
  ram matrix_c_8_14 (
    .addr0(c_addr_muxed_8_14_reg),
    .d0(c_data_8_14),
    .we0(we_c),
    .q0(data_from_out_mat_8_14),
    .clk(clk));

  //  BRAM matrix C8_15
  ram matrix_c_8_15 (
    .addr0(c_addr_muxed_8_15_reg),
    .d0(c_data_8_15),
    .we0(we_c),
    .q0(data_from_out_mat_8_15),
    .clk(clk));

  //  BRAM matrix C9_0
  ram matrix_c_9_0 (
    .addr0(c_addr_muxed_9_0_reg),
    .d0(c_data_9_0),
    .we0(we_c),
    .q0(data_from_out_mat_9_0),
    .clk(clk));

  //  BRAM matrix C9_1
  ram matrix_c_9_1 (
    .addr0(c_addr_muxed_9_1_reg),
    .d0(c_data_9_1),
    .we0(we_c),
    .q0(data_from_out_mat_9_1),
    .clk(clk));

  //  BRAM matrix C9_2
  ram matrix_c_9_2 (
    .addr0(c_addr_muxed_9_2_reg),
    .d0(c_data_9_2),
    .we0(we_c),
    .q0(data_from_out_mat_9_2),
    .clk(clk));

  //  BRAM matrix C9_3
  ram matrix_c_9_3 (
    .addr0(c_addr_muxed_9_3_reg),
    .d0(c_data_9_3),
    .we0(we_c),
    .q0(data_from_out_mat_9_3),
    .clk(clk));

  //  BRAM matrix C9_4
  ram matrix_c_9_4 (
    .addr0(c_addr_muxed_9_4_reg),
    .d0(c_data_9_4),
    .we0(we_c),
    .q0(data_from_out_mat_9_4),
    .clk(clk));

  //  BRAM matrix C9_5
  ram matrix_c_9_5 (
    .addr0(c_addr_muxed_9_5_reg),
    .d0(c_data_9_5),
    .we0(we_c),
    .q0(data_from_out_mat_9_5),
    .clk(clk));

  //  BRAM matrix C9_6
  ram matrix_c_9_6 (
    .addr0(c_addr_muxed_9_6_reg),
    .d0(c_data_9_6),
    .we0(we_c),
    .q0(data_from_out_mat_9_6),
    .clk(clk));

  //  BRAM matrix C9_7
  ram matrix_c_9_7 (
    .addr0(c_addr_muxed_9_7_reg),
    .d0(c_data_9_7),
    .we0(we_c),
    .q0(data_from_out_mat_9_7),
    .clk(clk));

  //  BRAM matrix C9_8
  ram matrix_c_9_8 (
    .addr0(c_addr_muxed_9_8_reg),
    .d0(c_data_9_8),
    .we0(we_c),
    .q0(data_from_out_mat_9_8),
    .clk(clk));

  //  BRAM matrix C9_9
  ram matrix_c_9_9 (
    .addr0(c_addr_muxed_9_9_reg),
    .d0(c_data_9_9),
    .we0(we_c),
    .q0(data_from_out_mat_9_9),
    .clk(clk));

  //  BRAM matrix C9_10
  ram matrix_c_9_10 (
    .addr0(c_addr_muxed_9_10_reg),
    .d0(c_data_9_10),
    .we0(we_c),
    .q0(data_from_out_mat_9_10),
    .clk(clk));

  //  BRAM matrix C9_11
  ram matrix_c_9_11 (
    .addr0(c_addr_muxed_9_11_reg),
    .d0(c_data_9_11),
    .we0(we_c),
    .q0(data_from_out_mat_9_11),
    .clk(clk));

  //  BRAM matrix C9_12
  ram matrix_c_9_12 (
    .addr0(c_addr_muxed_9_12_reg),
    .d0(c_data_9_12),
    .we0(we_c),
    .q0(data_from_out_mat_9_12),
    .clk(clk));

  //  BRAM matrix C9_13
  ram matrix_c_9_13 (
    .addr0(c_addr_muxed_9_13_reg),
    .d0(c_data_9_13),
    .we0(we_c),
    .q0(data_from_out_mat_9_13),
    .clk(clk));

  //  BRAM matrix C9_14
  ram matrix_c_9_14 (
    .addr0(c_addr_muxed_9_14_reg),
    .d0(c_data_9_14),
    .we0(we_c),
    .q0(data_from_out_mat_9_14),
    .clk(clk));

  //  BRAM matrix C9_15
  ram matrix_c_9_15 (
    .addr0(c_addr_muxed_9_15_reg),
    .d0(c_data_9_15),
    .we0(we_c),
    .q0(data_from_out_mat_9_15),
    .clk(clk));

  //  BRAM matrix C10_0
  ram matrix_c_10_0 (
    .addr0(c_addr_muxed_10_0_reg),
    .d0(c_data_10_0),
    .we0(we_c),
    .q0(data_from_out_mat_10_0),
    .clk(clk));

  //  BRAM matrix C10_1
  ram matrix_c_10_1 (
    .addr0(c_addr_muxed_10_1_reg),
    .d0(c_data_10_1),
    .we0(we_c),
    .q0(data_from_out_mat_10_1),
    .clk(clk));

  //  BRAM matrix C10_2
  ram matrix_c_10_2 (
    .addr0(c_addr_muxed_10_2_reg),
    .d0(c_data_10_2),
    .we0(we_c),
    .q0(data_from_out_mat_10_2),
    .clk(clk));

  //  BRAM matrix C10_3
  ram matrix_c_10_3 (
    .addr0(c_addr_muxed_10_3_reg),
    .d0(c_data_10_3),
    .we0(we_c),
    .q0(data_from_out_mat_10_3),
    .clk(clk));

  //  BRAM matrix C10_4
  ram matrix_c_10_4 (
    .addr0(c_addr_muxed_10_4_reg),
    .d0(c_data_10_4),
    .we0(we_c),
    .q0(data_from_out_mat_10_4),
    .clk(clk));

  //  BRAM matrix C10_5
  ram matrix_c_10_5 (
    .addr0(c_addr_muxed_10_5_reg),
    .d0(c_data_10_5),
    .we0(we_c),
    .q0(data_from_out_mat_10_5),
    .clk(clk));

  //  BRAM matrix C10_6
  ram matrix_c_10_6 (
    .addr0(c_addr_muxed_10_6_reg),
    .d0(c_data_10_6),
    .we0(we_c),
    .q0(data_from_out_mat_10_6),
    .clk(clk));

  //  BRAM matrix C10_7
  ram matrix_c_10_7 (
    .addr0(c_addr_muxed_10_7_reg),
    .d0(c_data_10_7),
    .we0(we_c),
    .q0(data_from_out_mat_10_7),
    .clk(clk));

  //  BRAM matrix C10_8
  ram matrix_c_10_8 (
    .addr0(c_addr_muxed_10_8_reg),
    .d0(c_data_10_8),
    .we0(we_c),
    .q0(data_from_out_mat_10_8),
    .clk(clk));

  //  BRAM matrix C10_9
  ram matrix_c_10_9 (
    .addr0(c_addr_muxed_10_9_reg),
    .d0(c_data_10_9),
    .we0(we_c),
    .q0(data_from_out_mat_10_9),
    .clk(clk));

  //  BRAM matrix C10_10
  ram matrix_c_10_10 (
    .addr0(c_addr_muxed_10_10_reg),
    .d0(c_data_10_10),
    .we0(we_c),
    .q0(data_from_out_mat_10_10),
    .clk(clk));

  //  BRAM matrix C10_11
  ram matrix_c_10_11 (
    .addr0(c_addr_muxed_10_11_reg),
    .d0(c_data_10_11),
    .we0(we_c),
    .q0(data_from_out_mat_10_11),
    .clk(clk));

  //  BRAM matrix C10_12
  ram matrix_c_10_12 (
    .addr0(c_addr_muxed_10_12_reg),
    .d0(c_data_10_12),
    .we0(we_c),
    .q0(data_from_out_mat_10_12),
    .clk(clk));

  //  BRAM matrix C10_13
  ram matrix_c_10_13 (
    .addr0(c_addr_muxed_10_13_reg),
    .d0(c_data_10_13),
    .we0(we_c),
    .q0(data_from_out_mat_10_13),
    .clk(clk));

  //  BRAM matrix C10_14
  ram matrix_c_10_14 (
    .addr0(c_addr_muxed_10_14_reg),
    .d0(c_data_10_14),
    .we0(we_c),
    .q0(data_from_out_mat_10_14),
    .clk(clk));

  //  BRAM matrix C10_15
  ram matrix_c_10_15 (
    .addr0(c_addr_muxed_10_15_reg),
    .d0(c_data_10_15),
    .we0(we_c),
    .q0(data_from_out_mat_10_15),
    .clk(clk));

  //  BRAM matrix C11_0
  ram matrix_c_11_0 (
    .addr0(c_addr_muxed_11_0_reg),
    .d0(c_data_11_0),
    .we0(we_c),
    .q0(data_from_out_mat_11_0),
    .clk(clk));

  //  BRAM matrix C11_1
  ram matrix_c_11_1 (
    .addr0(c_addr_muxed_11_1_reg),
    .d0(c_data_11_1),
    .we0(we_c),
    .q0(data_from_out_mat_11_1),
    .clk(clk));

  //  BRAM matrix C11_2
  ram matrix_c_11_2 (
    .addr0(c_addr_muxed_11_2_reg),
    .d0(c_data_11_2),
    .we0(we_c),
    .q0(data_from_out_mat_11_2),
    .clk(clk));

  //  BRAM matrix C11_3
  ram matrix_c_11_3 (
    .addr0(c_addr_muxed_11_3_reg),
    .d0(c_data_11_3),
    .we0(we_c),
    .q0(data_from_out_mat_11_3),
    .clk(clk));

  //  BRAM matrix C11_4
  ram matrix_c_11_4 (
    .addr0(c_addr_muxed_11_4_reg),
    .d0(c_data_11_4),
    .we0(we_c),
    .q0(data_from_out_mat_11_4),
    .clk(clk));

  //  BRAM matrix C11_5
  ram matrix_c_11_5 (
    .addr0(c_addr_muxed_11_5_reg),
    .d0(c_data_11_5),
    .we0(we_c),
    .q0(data_from_out_mat_11_5),
    .clk(clk));

  //  BRAM matrix C11_6
  ram matrix_c_11_6 (
    .addr0(c_addr_muxed_11_6_reg),
    .d0(c_data_11_6),
    .we0(we_c),
    .q0(data_from_out_mat_11_6),
    .clk(clk));

  //  BRAM matrix C11_7
  ram matrix_c_11_7 (
    .addr0(c_addr_muxed_11_7_reg),
    .d0(c_data_11_7),
    .we0(we_c),
    .q0(data_from_out_mat_11_7),
    .clk(clk));

  //  BRAM matrix C11_8
  ram matrix_c_11_8 (
    .addr0(c_addr_muxed_11_8_reg),
    .d0(c_data_11_8),
    .we0(we_c),
    .q0(data_from_out_mat_11_8),
    .clk(clk));

  //  BRAM matrix C11_9
  ram matrix_c_11_9 (
    .addr0(c_addr_muxed_11_9_reg),
    .d0(c_data_11_9),
    .we0(we_c),
    .q0(data_from_out_mat_11_9),
    .clk(clk));

  //  BRAM matrix C11_10
  ram matrix_c_11_10 (
    .addr0(c_addr_muxed_11_10_reg),
    .d0(c_data_11_10),
    .we0(we_c),
    .q0(data_from_out_mat_11_10),
    .clk(clk));

  //  BRAM matrix C11_11
  ram matrix_c_11_11 (
    .addr0(c_addr_muxed_11_11_reg),
    .d0(c_data_11_11),
    .we0(we_c),
    .q0(data_from_out_mat_11_11),
    .clk(clk));

  //  BRAM matrix C11_12
  ram matrix_c_11_12 (
    .addr0(c_addr_muxed_11_12_reg),
    .d0(c_data_11_12),
    .we0(we_c),
    .q0(data_from_out_mat_11_12),
    .clk(clk));

  //  BRAM matrix C11_13
  ram matrix_c_11_13 (
    .addr0(c_addr_muxed_11_13_reg),
    .d0(c_data_11_13),
    .we0(we_c),
    .q0(data_from_out_mat_11_13),
    .clk(clk));

  //  BRAM matrix C11_14
  ram matrix_c_11_14 (
    .addr0(c_addr_muxed_11_14_reg),
    .d0(c_data_11_14),
    .we0(we_c),
    .q0(data_from_out_mat_11_14),
    .clk(clk));

  //  BRAM matrix C11_15
  ram matrix_c_11_15 (
    .addr0(c_addr_muxed_11_15_reg),
    .d0(c_data_11_15),
    .we0(we_c),
    .q0(data_from_out_mat_11_15),
    .clk(clk));

  //  BRAM matrix C12_0
  ram matrix_c_12_0 (
    .addr0(c_addr_muxed_12_0_reg),
    .d0(c_data_12_0),
    .we0(we_c),
    .q0(data_from_out_mat_12_0),
    .clk(clk));

  //  BRAM matrix C12_1
  ram matrix_c_12_1 (
    .addr0(c_addr_muxed_12_1_reg),
    .d0(c_data_12_1),
    .we0(we_c),
    .q0(data_from_out_mat_12_1),
    .clk(clk));

  //  BRAM matrix C12_2
  ram matrix_c_12_2 (
    .addr0(c_addr_muxed_12_2_reg),
    .d0(c_data_12_2),
    .we0(we_c),
    .q0(data_from_out_mat_12_2),
    .clk(clk));

  //  BRAM matrix C12_3
  ram matrix_c_12_3 (
    .addr0(c_addr_muxed_12_3_reg),
    .d0(c_data_12_3),
    .we0(we_c),
    .q0(data_from_out_mat_12_3),
    .clk(clk));

  //  BRAM matrix C12_4
  ram matrix_c_12_4 (
    .addr0(c_addr_muxed_12_4_reg),
    .d0(c_data_12_4),
    .we0(we_c),
    .q0(data_from_out_mat_12_4),
    .clk(clk));

  //  BRAM matrix C12_5
  ram matrix_c_12_5 (
    .addr0(c_addr_muxed_12_5_reg),
    .d0(c_data_12_5),
    .we0(we_c),
    .q0(data_from_out_mat_12_5),
    .clk(clk));

  //  BRAM matrix C12_6
  ram matrix_c_12_6 (
    .addr0(c_addr_muxed_12_6_reg),
    .d0(c_data_12_6),
    .we0(we_c),
    .q0(data_from_out_mat_12_6),
    .clk(clk));

  //  BRAM matrix C12_7
  ram matrix_c_12_7 (
    .addr0(c_addr_muxed_12_7_reg),
    .d0(c_data_12_7),
    .we0(we_c),
    .q0(data_from_out_mat_12_7),
    .clk(clk));

  //  BRAM matrix C12_8
  ram matrix_c_12_8 (
    .addr0(c_addr_muxed_12_8_reg),
    .d0(c_data_12_8),
    .we0(we_c),
    .q0(data_from_out_mat_12_8),
    .clk(clk));

  //  BRAM matrix C12_9
  ram matrix_c_12_9 (
    .addr0(c_addr_muxed_12_9_reg),
    .d0(c_data_12_9),
    .we0(we_c),
    .q0(data_from_out_mat_12_9),
    .clk(clk));

  //  BRAM matrix C12_10
  ram matrix_c_12_10 (
    .addr0(c_addr_muxed_12_10_reg),
    .d0(c_data_12_10),
    .we0(we_c),
    .q0(data_from_out_mat_12_10),
    .clk(clk));

  //  BRAM matrix C12_11
  ram matrix_c_12_11 (
    .addr0(c_addr_muxed_12_11_reg),
    .d0(c_data_12_11),
    .we0(we_c),
    .q0(data_from_out_mat_12_11),
    .clk(clk));

  //  BRAM matrix C12_12
  ram matrix_c_12_12 (
    .addr0(c_addr_muxed_12_12_reg),
    .d0(c_data_12_12),
    .we0(we_c),
    .q0(data_from_out_mat_12_12),
    .clk(clk));

  //  BRAM matrix C12_13
  ram matrix_c_12_13 (
    .addr0(c_addr_muxed_12_13_reg),
    .d0(c_data_12_13),
    .we0(we_c),
    .q0(data_from_out_mat_12_13),
    .clk(clk));

  //  BRAM matrix C12_14
  ram matrix_c_12_14 (
    .addr0(c_addr_muxed_12_14_reg),
    .d0(c_data_12_14),
    .we0(we_c),
    .q0(data_from_out_mat_12_14),
    .clk(clk));

  //  BRAM matrix C12_15
  ram matrix_c_12_15 (
    .addr0(c_addr_muxed_12_15_reg),
    .d0(c_data_12_15),
    .we0(we_c),
    .q0(data_from_out_mat_12_15),
    .clk(clk));

  //  BRAM matrix C13_0
  ram matrix_c_13_0 (
    .addr0(c_addr_muxed_13_0_reg),
    .d0(c_data_13_0),
    .we0(we_c),
    .q0(data_from_out_mat_13_0),
    .clk(clk));

  //  BRAM matrix C13_1
  ram matrix_c_13_1 (
    .addr0(c_addr_muxed_13_1_reg),
    .d0(c_data_13_1),
    .we0(we_c),
    .q0(data_from_out_mat_13_1),
    .clk(clk));

  //  BRAM matrix C13_2
  ram matrix_c_13_2 (
    .addr0(c_addr_muxed_13_2_reg),
    .d0(c_data_13_2),
    .we0(we_c),
    .q0(data_from_out_mat_13_2),
    .clk(clk));

  //  BRAM matrix C13_3
  ram matrix_c_13_3 (
    .addr0(c_addr_muxed_13_3_reg),
    .d0(c_data_13_3),
    .we0(we_c),
    .q0(data_from_out_mat_13_3),
    .clk(clk));

  //  BRAM matrix C13_4
  ram matrix_c_13_4 (
    .addr0(c_addr_muxed_13_4_reg),
    .d0(c_data_13_4),
    .we0(we_c),
    .q0(data_from_out_mat_13_4),
    .clk(clk));

  //  BRAM matrix C13_5
  ram matrix_c_13_5 (
    .addr0(c_addr_muxed_13_5_reg),
    .d0(c_data_13_5),
    .we0(we_c),
    .q0(data_from_out_mat_13_5),
    .clk(clk));

  //  BRAM matrix C13_6
  ram matrix_c_13_6 (
    .addr0(c_addr_muxed_13_6_reg),
    .d0(c_data_13_6),
    .we0(we_c),
    .q0(data_from_out_mat_13_6),
    .clk(clk));

  //  BRAM matrix C13_7
  ram matrix_c_13_7 (
    .addr0(c_addr_muxed_13_7_reg),
    .d0(c_data_13_7),
    .we0(we_c),
    .q0(data_from_out_mat_13_7),
    .clk(clk));

  //  BRAM matrix C13_8
  ram matrix_c_13_8 (
    .addr0(c_addr_muxed_13_8_reg),
    .d0(c_data_13_8),
    .we0(we_c),
    .q0(data_from_out_mat_13_8),
    .clk(clk));

  //  BRAM matrix C13_9
  ram matrix_c_13_9 (
    .addr0(c_addr_muxed_13_9_reg),
    .d0(c_data_13_9),
    .we0(we_c),
    .q0(data_from_out_mat_13_9),
    .clk(clk));

  //  BRAM matrix C13_10
  ram matrix_c_13_10 (
    .addr0(c_addr_muxed_13_10_reg),
    .d0(c_data_13_10),
    .we0(we_c),
    .q0(data_from_out_mat_13_10),
    .clk(clk));

  //  BRAM matrix C13_11
  ram matrix_c_13_11 (
    .addr0(c_addr_muxed_13_11_reg),
    .d0(c_data_13_11),
    .we0(we_c),
    .q0(data_from_out_mat_13_11),
    .clk(clk));

  //  BRAM matrix C13_12
  ram matrix_c_13_12 (
    .addr0(c_addr_muxed_13_12_reg),
    .d0(c_data_13_12),
    .we0(we_c),
    .q0(data_from_out_mat_13_12),
    .clk(clk));

  //  BRAM matrix C13_13
  ram matrix_c_13_13 (
    .addr0(c_addr_muxed_13_13_reg),
    .d0(c_data_13_13),
    .we0(we_c),
    .q0(data_from_out_mat_13_13),
    .clk(clk));

  //  BRAM matrix C13_14
  ram matrix_c_13_14 (
    .addr0(c_addr_muxed_13_14_reg),
    .d0(c_data_13_14),
    .we0(we_c),
    .q0(data_from_out_mat_13_14),
    .clk(clk));

  //  BRAM matrix C13_15
  ram matrix_c_13_15 (
    .addr0(c_addr_muxed_13_15_reg),
    .d0(c_data_13_15),
    .we0(we_c),
    .q0(data_from_out_mat_13_15),
    .clk(clk));

  //  BRAM matrix C14_0
  ram matrix_c_14_0 (
    .addr0(c_addr_muxed_14_0_reg),
    .d0(c_data_14_0),
    .we0(we_c),
    .q0(data_from_out_mat_14_0),
    .clk(clk));

  //  BRAM matrix C14_1
  ram matrix_c_14_1 (
    .addr0(c_addr_muxed_14_1_reg),
    .d0(c_data_14_1),
    .we0(we_c),
    .q0(data_from_out_mat_14_1),
    .clk(clk));

  //  BRAM matrix C14_2
  ram matrix_c_14_2 (
    .addr0(c_addr_muxed_14_2_reg),
    .d0(c_data_14_2),
    .we0(we_c),
    .q0(data_from_out_mat_14_2),
    .clk(clk));

  //  BRAM matrix C14_3
  ram matrix_c_14_3 (
    .addr0(c_addr_muxed_14_3_reg),
    .d0(c_data_14_3),
    .we0(we_c),
    .q0(data_from_out_mat_14_3),
    .clk(clk));

  //  BRAM matrix C14_4
  ram matrix_c_14_4 (
    .addr0(c_addr_muxed_14_4_reg),
    .d0(c_data_14_4),
    .we0(we_c),
    .q0(data_from_out_mat_14_4),
    .clk(clk));

  //  BRAM matrix C14_5
  ram matrix_c_14_5 (
    .addr0(c_addr_muxed_14_5_reg),
    .d0(c_data_14_5),
    .we0(we_c),
    .q0(data_from_out_mat_14_5),
    .clk(clk));

  //  BRAM matrix C14_6
  ram matrix_c_14_6 (
    .addr0(c_addr_muxed_14_6_reg),
    .d0(c_data_14_6),
    .we0(we_c),
    .q0(data_from_out_mat_14_6),
    .clk(clk));

  //  BRAM matrix C14_7
  ram matrix_c_14_7 (
    .addr0(c_addr_muxed_14_7_reg),
    .d0(c_data_14_7),
    .we0(we_c),
    .q0(data_from_out_mat_14_7),
    .clk(clk));

  //  BRAM matrix C14_8
  ram matrix_c_14_8 (
    .addr0(c_addr_muxed_14_8_reg),
    .d0(c_data_14_8),
    .we0(we_c),
    .q0(data_from_out_mat_14_8),
    .clk(clk));

  //  BRAM matrix C14_9
  ram matrix_c_14_9 (
    .addr0(c_addr_muxed_14_9_reg),
    .d0(c_data_14_9),
    .we0(we_c),
    .q0(data_from_out_mat_14_9),
    .clk(clk));

  //  BRAM matrix C14_10
  ram matrix_c_14_10 (
    .addr0(c_addr_muxed_14_10_reg),
    .d0(c_data_14_10),
    .we0(we_c),
    .q0(data_from_out_mat_14_10),
    .clk(clk));

  //  BRAM matrix C14_11
  ram matrix_c_14_11 (
    .addr0(c_addr_muxed_14_11_reg),
    .d0(c_data_14_11),
    .we0(we_c),
    .q0(data_from_out_mat_14_11),
    .clk(clk));

  //  BRAM matrix C14_12
  ram matrix_c_14_12 (
    .addr0(c_addr_muxed_14_12_reg),
    .d0(c_data_14_12),
    .we0(we_c),
    .q0(data_from_out_mat_14_12),
    .clk(clk));

  //  BRAM matrix C14_13
  ram matrix_c_14_13 (
    .addr0(c_addr_muxed_14_13_reg),
    .d0(c_data_14_13),
    .we0(we_c),
    .q0(data_from_out_mat_14_13),
    .clk(clk));

  //  BRAM matrix C14_14
  ram matrix_c_14_14 (
    .addr0(c_addr_muxed_14_14_reg),
    .d0(c_data_14_14),
    .we0(we_c),
    .q0(data_from_out_mat_14_14),
    .clk(clk));

  //  BRAM matrix C14_15
  ram matrix_c_14_15 (
    .addr0(c_addr_muxed_14_15_reg),
    .d0(c_data_14_15),
    .we0(we_c),
    .q0(data_from_out_mat_14_15),
    .clk(clk));

  //  BRAM matrix C15_0
  ram matrix_c_15_0 (
    .addr0(c_addr_muxed_15_0_reg),
    .d0(c_data_15_0),
    .we0(we_c),
    .q0(data_from_out_mat_15_0),
    .clk(clk));

  //  BRAM matrix C15_1
  ram matrix_c_15_1 (
    .addr0(c_addr_muxed_15_1_reg),
    .d0(c_data_15_1),
    .we0(we_c),
    .q0(data_from_out_mat_15_1),
    .clk(clk));

  //  BRAM matrix C15_2
  ram matrix_c_15_2 (
    .addr0(c_addr_muxed_15_2_reg),
    .d0(c_data_15_2),
    .we0(we_c),
    .q0(data_from_out_mat_15_2),
    .clk(clk));

  //  BRAM matrix C15_3
  ram matrix_c_15_3 (
    .addr0(c_addr_muxed_15_3_reg),
    .d0(c_data_15_3),
    .we0(we_c),
    .q0(data_from_out_mat_15_3),
    .clk(clk));

  //  BRAM matrix C15_4
  ram matrix_c_15_4 (
    .addr0(c_addr_muxed_15_4_reg),
    .d0(c_data_15_4),
    .we0(we_c),
    .q0(data_from_out_mat_15_4),
    .clk(clk));

  //  BRAM matrix C15_5
  ram matrix_c_15_5 (
    .addr0(c_addr_muxed_15_5_reg),
    .d0(c_data_15_5),
    .we0(we_c),
    .q0(data_from_out_mat_15_5),
    .clk(clk));

  //  BRAM matrix C15_6
  ram matrix_c_15_6 (
    .addr0(c_addr_muxed_15_6_reg),
    .d0(c_data_15_6),
    .we0(we_c),
    .q0(data_from_out_mat_15_6),
    .clk(clk));

  //  BRAM matrix C15_7
  ram matrix_c_15_7 (
    .addr0(c_addr_muxed_15_7_reg),
    .d0(c_data_15_7),
    .we0(we_c),
    .q0(data_from_out_mat_15_7),
    .clk(clk));

  //  BRAM matrix C15_8
  ram matrix_c_15_8 (
    .addr0(c_addr_muxed_15_8_reg),
    .d0(c_data_15_8),
    .we0(we_c),
    .q0(data_from_out_mat_15_8),
    .clk(clk));

  //  BRAM matrix C15_9
  ram matrix_c_15_9 (
    .addr0(c_addr_muxed_15_9_reg),
    .d0(c_data_15_9),
    .we0(we_c),
    .q0(data_from_out_mat_15_9),
    .clk(clk));

  //  BRAM matrix C15_10
  ram matrix_c_15_10 (
    .addr0(c_addr_muxed_15_10_reg),
    .d0(c_data_15_10),
    .we0(we_c),
    .q0(data_from_out_mat_15_10),
    .clk(clk));

  //  BRAM matrix C15_11
  ram matrix_c_15_11 (
    .addr0(c_addr_muxed_15_11_reg),
    .d0(c_data_15_11),
    .we0(we_c),
    .q0(data_from_out_mat_15_11),
    .clk(clk));

  //  BRAM matrix C15_12
  ram matrix_c_15_12 (
    .addr0(c_addr_muxed_15_12_reg),
    .d0(c_data_15_12),
    .we0(we_c),
    .q0(data_from_out_mat_15_12),
    .clk(clk));

  //  BRAM matrix C15_13
  ram matrix_c_15_13 (
    .addr0(c_addr_muxed_15_13_reg),
    .d0(c_data_15_13),
    .we0(we_c),
    .q0(data_from_out_mat_15_13),
    .clk(clk));

  //  BRAM matrix C15_14
  ram matrix_c_15_14 (
    .addr0(c_addr_muxed_15_14_reg),
    .d0(c_data_15_14),
    .we0(we_c),
    .q0(data_from_out_mat_15_14),
    .clk(clk));

  //  BRAM matrix C15_15
  ram matrix_c_15_15 (
    .addr0(c_addr_muxed_15_15_reg),
    .d0(c_data_15_15),
    .we0(we_c),
    .q0(data_from_out_mat_15_15),
    .clk(clk));

/////////////////////////////////////////////////
// The 64x64 matmul instantiation
/////////////////////////////////////////////////

matmul_64x64_systolic u_matmul_64x64_systolic (
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul),
  .a_data_0_0(a_data_0_0),
  .a_addr_0_0(a_addr_0_0),
  .b_data_0_0(b_data_0_0),
  .b_addr_0_0(b_addr_0_0),
  .a_data_1_0(a_data_1_0),
  .a_addr_1_0(a_addr_1_0),
  .b_data_0_1(b_data_0_1),
  .b_addr_0_1(b_addr_0_1),
  .a_data_2_0(a_data_2_0),
  .a_addr_2_0(a_addr_2_0),
  .b_data_0_2(b_data_0_2),
  .b_addr_0_2(b_addr_0_2),
  .a_data_3_0(a_data_3_0),
  .a_addr_3_0(a_addr_3_0),
  .b_data_0_3(b_data_0_3),
  .b_addr_0_3(b_addr_0_3),
  .a_data_4_0(a_data_4_0),
  .a_addr_4_0(a_addr_4_0),
  .b_data_0_4(b_data_0_4),
  .b_addr_0_4(b_addr_0_4),
  .a_data_5_0(a_data_5_0),
  .a_addr_5_0(a_addr_5_0),
  .b_data_0_5(b_data_0_5),
  .b_addr_0_5(b_addr_0_5),
  .a_data_6_0(a_data_6_0),
  .a_addr_6_0(a_addr_6_0),
  .b_data_0_6(b_data_0_6),
  .b_addr_0_6(b_addr_0_6),
  .a_data_7_0(a_data_7_0),
  .a_addr_7_0(a_addr_7_0),
  .b_data_0_7(b_data_0_7),
  .b_addr_0_7(b_addr_0_7),
  .a_data_8_0(a_data_8_0),
  .a_addr_8_0(a_addr_8_0),
  .b_data_0_8(b_data_0_8),
  .b_addr_0_8(b_addr_0_8),
  .a_data_9_0(a_data_9_0),
  .a_addr_9_0(a_addr_9_0),
  .b_data_0_9(b_data_0_9),
  .b_addr_0_9(b_addr_0_9),
  .a_data_10_0(a_data_10_0),
  .a_addr_10_0(a_addr_10_0),
  .b_data_0_10(b_data_0_10),
  .b_addr_0_10(b_addr_0_10),
  .a_data_11_0(a_data_11_0),
  .a_addr_11_0(a_addr_11_0),
  .b_data_0_11(b_data_0_11),
  .b_addr_0_11(b_addr_0_11),
  .a_data_12_0(a_data_12_0),
  .a_addr_12_0(a_addr_12_0),
  .b_data_0_12(b_data_0_12),
  .b_addr_0_12(b_addr_0_12),
  .a_data_13_0(a_data_13_0),
  .a_addr_13_0(a_addr_13_0),
  .b_data_0_13(b_data_0_13),
  .b_addr_0_13(b_addr_0_13),
  .a_data_14_0(a_data_14_0),
  .a_addr_14_0(a_addr_14_0),
  .b_data_0_14(b_data_0_14),
  .b_addr_0_14(b_addr_0_14),
  .a_data_15_0(a_data_15_0),
  .a_addr_15_0(a_addr_15_0),
  .b_data_0_15(b_data_0_15),
  .b_addr_0_15(b_addr_0_15),

  .c_data_0_0(c_data_0_0),
  .c_addr_0_0(c_addr_0_0),
  .c_data_0_1(c_data_0_1),
  .c_addr_0_1(c_addr_0_1),
  .c_data_0_2(c_data_0_2),
  .c_addr_0_2(c_addr_0_2),
  .c_data_0_3(c_data_0_3),
  .c_addr_0_3(c_addr_0_3),
  .c_data_0_4(c_data_0_4),
  .c_addr_0_4(c_addr_0_4),
  .c_data_0_5(c_data_0_5),
  .c_addr_0_5(c_addr_0_5),
  .c_data_0_6(c_data_0_6),
  .c_addr_0_6(c_addr_0_6),
  .c_data_0_7(c_data_0_7),
  .c_addr_0_7(c_addr_0_7),
  .c_data_0_8(c_data_0_8),
  .c_addr_0_8(c_addr_0_8),
  .c_data_0_9(c_data_0_9),
  .c_addr_0_9(c_addr_0_9),
  .c_data_0_10(c_data_0_10),
  .c_addr_0_10(c_addr_0_10),
  .c_data_0_11(c_data_0_11),
  .c_addr_0_11(c_addr_0_11),
  .c_data_0_12(c_data_0_12),
  .c_addr_0_12(c_addr_0_12),
  .c_data_0_13(c_data_0_13),
  .c_addr_0_13(c_addr_0_13),
  .c_data_0_14(c_data_0_14),
  .c_addr_0_14(c_addr_0_14),
  .c_data_0_15(c_data_0_15),
  .c_addr_0_15(c_addr_0_15),
  .c_data_1_0(c_data_1_0),
  .c_addr_1_0(c_addr_1_0),
  .c_data_1_1(c_data_1_1),
  .c_addr_1_1(c_addr_1_1),
  .c_data_1_2(c_data_1_2),
  .c_addr_1_2(c_addr_1_2),
  .c_data_1_3(c_data_1_3),
  .c_addr_1_3(c_addr_1_3),
  .c_data_1_4(c_data_1_4),
  .c_addr_1_4(c_addr_1_4),
  .c_data_1_5(c_data_1_5),
  .c_addr_1_5(c_addr_1_5),
  .c_data_1_6(c_data_1_6),
  .c_addr_1_6(c_addr_1_6),
  .c_data_1_7(c_data_1_7),
  .c_addr_1_7(c_addr_1_7),
  .c_data_1_8(c_data_1_8),
  .c_addr_1_8(c_addr_1_8),
  .c_data_1_9(c_data_1_9),
  .c_addr_1_9(c_addr_1_9),
  .c_data_1_10(c_data_1_10),
  .c_addr_1_10(c_addr_1_10),
  .c_data_1_11(c_data_1_11),
  .c_addr_1_11(c_addr_1_11),
  .c_data_1_12(c_data_1_12),
  .c_addr_1_12(c_addr_1_12),
  .c_data_1_13(c_data_1_13),
  .c_addr_1_13(c_addr_1_13),
  .c_data_1_14(c_data_1_14),
  .c_addr_1_14(c_addr_1_14),
  .c_data_1_15(c_data_1_15),
  .c_addr_1_15(c_addr_1_15),
  .c_data_2_0(c_data_2_0),
  .c_addr_2_0(c_addr_2_0),
  .c_data_2_1(c_data_2_1),
  .c_addr_2_1(c_addr_2_1),
  .c_data_2_2(c_data_2_2),
  .c_addr_2_2(c_addr_2_2),
  .c_data_2_3(c_data_2_3),
  .c_addr_2_3(c_addr_2_3),
  .c_data_2_4(c_data_2_4),
  .c_addr_2_4(c_addr_2_4),
  .c_data_2_5(c_data_2_5),
  .c_addr_2_5(c_addr_2_5),
  .c_data_2_6(c_data_2_6),
  .c_addr_2_6(c_addr_2_6),
  .c_data_2_7(c_data_2_7),
  .c_addr_2_7(c_addr_2_7),
  .c_data_2_8(c_data_2_8),
  .c_addr_2_8(c_addr_2_8),
  .c_data_2_9(c_data_2_9),
  .c_addr_2_9(c_addr_2_9),
  .c_data_2_10(c_data_2_10),
  .c_addr_2_10(c_addr_2_10),
  .c_data_2_11(c_data_2_11),
  .c_addr_2_11(c_addr_2_11),
  .c_data_2_12(c_data_2_12),
  .c_addr_2_12(c_addr_2_12),
  .c_data_2_13(c_data_2_13),
  .c_addr_2_13(c_addr_2_13),
  .c_data_2_14(c_data_2_14),
  .c_addr_2_14(c_addr_2_14),
  .c_data_2_15(c_data_2_15),
  .c_addr_2_15(c_addr_2_15),
  .c_data_3_0(c_data_3_0),
  .c_addr_3_0(c_addr_3_0),
  .c_data_3_1(c_data_3_1),
  .c_addr_3_1(c_addr_3_1),
  .c_data_3_2(c_data_3_2),
  .c_addr_3_2(c_addr_3_2),
  .c_data_3_3(c_data_3_3),
  .c_addr_3_3(c_addr_3_3),
  .c_data_3_4(c_data_3_4),
  .c_addr_3_4(c_addr_3_4),
  .c_data_3_5(c_data_3_5),
  .c_addr_3_5(c_addr_3_5),
  .c_data_3_6(c_data_3_6),
  .c_addr_3_6(c_addr_3_6),
  .c_data_3_7(c_data_3_7),
  .c_addr_3_7(c_addr_3_7),
  .c_data_3_8(c_data_3_8),
  .c_addr_3_8(c_addr_3_8),
  .c_data_3_9(c_data_3_9),
  .c_addr_3_9(c_addr_3_9),
  .c_data_3_10(c_data_3_10),
  .c_addr_3_10(c_addr_3_10),
  .c_data_3_11(c_data_3_11),
  .c_addr_3_11(c_addr_3_11),
  .c_data_3_12(c_data_3_12),
  .c_addr_3_12(c_addr_3_12),
  .c_data_3_13(c_data_3_13),
  .c_addr_3_13(c_addr_3_13),
  .c_data_3_14(c_data_3_14),
  .c_addr_3_14(c_addr_3_14),
  .c_data_3_15(c_data_3_15),
  .c_addr_3_15(c_addr_3_15),
  .c_data_4_0(c_data_4_0),
  .c_addr_4_0(c_addr_4_0),
  .c_data_4_1(c_data_4_1),
  .c_addr_4_1(c_addr_4_1),
  .c_data_4_2(c_data_4_2),
  .c_addr_4_2(c_addr_4_2),
  .c_data_4_3(c_data_4_3),
  .c_addr_4_3(c_addr_4_3),
  .c_data_4_4(c_data_4_4),
  .c_addr_4_4(c_addr_4_4),
  .c_data_4_5(c_data_4_5),
  .c_addr_4_5(c_addr_4_5),
  .c_data_4_6(c_data_4_6),
  .c_addr_4_6(c_addr_4_6),
  .c_data_4_7(c_data_4_7),
  .c_addr_4_7(c_addr_4_7),
  .c_data_4_8(c_data_4_8),
  .c_addr_4_8(c_addr_4_8),
  .c_data_4_9(c_data_4_9),
  .c_addr_4_9(c_addr_4_9),
  .c_data_4_10(c_data_4_10),
  .c_addr_4_10(c_addr_4_10),
  .c_data_4_11(c_data_4_11),
  .c_addr_4_11(c_addr_4_11),
  .c_data_4_12(c_data_4_12),
  .c_addr_4_12(c_addr_4_12),
  .c_data_4_13(c_data_4_13),
  .c_addr_4_13(c_addr_4_13),
  .c_data_4_14(c_data_4_14),
  .c_addr_4_14(c_addr_4_14),
  .c_data_4_15(c_data_4_15),
  .c_addr_4_15(c_addr_4_15),
  .c_data_5_0(c_data_5_0),
  .c_addr_5_0(c_addr_5_0),
  .c_data_5_1(c_data_5_1),
  .c_addr_5_1(c_addr_5_1),
  .c_data_5_2(c_data_5_2),
  .c_addr_5_2(c_addr_5_2),
  .c_data_5_3(c_data_5_3),
  .c_addr_5_3(c_addr_5_3),
  .c_data_5_4(c_data_5_4),
  .c_addr_5_4(c_addr_5_4),
  .c_data_5_5(c_data_5_5),
  .c_addr_5_5(c_addr_5_5),
  .c_data_5_6(c_data_5_6),
  .c_addr_5_6(c_addr_5_6),
  .c_data_5_7(c_data_5_7),
  .c_addr_5_7(c_addr_5_7),
  .c_data_5_8(c_data_5_8),
  .c_addr_5_8(c_addr_5_8),
  .c_data_5_9(c_data_5_9),
  .c_addr_5_9(c_addr_5_9),
  .c_data_5_10(c_data_5_10),
  .c_addr_5_10(c_addr_5_10),
  .c_data_5_11(c_data_5_11),
  .c_addr_5_11(c_addr_5_11),
  .c_data_5_12(c_data_5_12),
  .c_addr_5_12(c_addr_5_12),
  .c_data_5_13(c_data_5_13),
  .c_addr_5_13(c_addr_5_13),
  .c_data_5_14(c_data_5_14),
  .c_addr_5_14(c_addr_5_14),
  .c_data_5_15(c_data_5_15),
  .c_addr_5_15(c_addr_5_15),
  .c_data_6_0(c_data_6_0),
  .c_addr_6_0(c_addr_6_0),
  .c_data_6_1(c_data_6_1),
  .c_addr_6_1(c_addr_6_1),
  .c_data_6_2(c_data_6_2),
  .c_addr_6_2(c_addr_6_2),
  .c_data_6_3(c_data_6_3),
  .c_addr_6_3(c_addr_6_3),
  .c_data_6_4(c_data_6_4),
  .c_addr_6_4(c_addr_6_4),
  .c_data_6_5(c_data_6_5),
  .c_addr_6_5(c_addr_6_5),
  .c_data_6_6(c_data_6_6),
  .c_addr_6_6(c_addr_6_6),
  .c_data_6_7(c_data_6_7),
  .c_addr_6_7(c_addr_6_7),
  .c_data_6_8(c_data_6_8),
  .c_addr_6_8(c_addr_6_8),
  .c_data_6_9(c_data_6_9),
  .c_addr_6_9(c_addr_6_9),
  .c_data_6_10(c_data_6_10),
  .c_addr_6_10(c_addr_6_10),
  .c_data_6_11(c_data_6_11),
  .c_addr_6_11(c_addr_6_11),
  .c_data_6_12(c_data_6_12),
  .c_addr_6_12(c_addr_6_12),
  .c_data_6_13(c_data_6_13),
  .c_addr_6_13(c_addr_6_13),
  .c_data_6_14(c_data_6_14),
  .c_addr_6_14(c_addr_6_14),
  .c_data_6_15(c_data_6_15),
  .c_addr_6_15(c_addr_6_15),
  .c_data_7_0(c_data_7_0),
  .c_addr_7_0(c_addr_7_0),
  .c_data_7_1(c_data_7_1),
  .c_addr_7_1(c_addr_7_1),
  .c_data_7_2(c_data_7_2),
  .c_addr_7_2(c_addr_7_2),
  .c_data_7_3(c_data_7_3),
  .c_addr_7_3(c_addr_7_3),
  .c_data_7_4(c_data_7_4),
  .c_addr_7_4(c_addr_7_4),
  .c_data_7_5(c_data_7_5),
  .c_addr_7_5(c_addr_7_5),
  .c_data_7_6(c_data_7_6),
  .c_addr_7_6(c_addr_7_6),
  .c_data_7_7(c_data_7_7),
  .c_addr_7_7(c_addr_7_7),
  .c_data_7_8(c_data_7_8),
  .c_addr_7_8(c_addr_7_8),
  .c_data_7_9(c_data_7_9),
  .c_addr_7_9(c_addr_7_9),
  .c_data_7_10(c_data_7_10),
  .c_addr_7_10(c_addr_7_10),
  .c_data_7_11(c_data_7_11),
  .c_addr_7_11(c_addr_7_11),
  .c_data_7_12(c_data_7_12),
  .c_addr_7_12(c_addr_7_12),
  .c_data_7_13(c_data_7_13),
  .c_addr_7_13(c_addr_7_13),
  .c_data_7_14(c_data_7_14),
  .c_addr_7_14(c_addr_7_14),
  .c_data_7_15(c_data_7_15),
  .c_addr_7_15(c_addr_7_15),
  .c_data_8_0(c_data_8_0),
  .c_addr_8_0(c_addr_8_0),
  .c_data_8_1(c_data_8_1),
  .c_addr_8_1(c_addr_8_1),
  .c_data_8_2(c_data_8_2),
  .c_addr_8_2(c_addr_8_2),
  .c_data_8_3(c_data_8_3),
  .c_addr_8_3(c_addr_8_3),
  .c_data_8_4(c_data_8_4),
  .c_addr_8_4(c_addr_8_4),
  .c_data_8_5(c_data_8_5),
  .c_addr_8_5(c_addr_8_5),
  .c_data_8_6(c_data_8_6),
  .c_addr_8_6(c_addr_8_6),
  .c_data_8_7(c_data_8_7),
  .c_addr_8_7(c_addr_8_7),
  .c_data_8_8(c_data_8_8),
  .c_addr_8_8(c_addr_8_8),
  .c_data_8_9(c_data_8_9),
  .c_addr_8_9(c_addr_8_9),
  .c_data_8_10(c_data_8_10),
  .c_addr_8_10(c_addr_8_10),
  .c_data_8_11(c_data_8_11),
  .c_addr_8_11(c_addr_8_11),
  .c_data_8_12(c_data_8_12),
  .c_addr_8_12(c_addr_8_12),
  .c_data_8_13(c_data_8_13),
  .c_addr_8_13(c_addr_8_13),
  .c_data_8_14(c_data_8_14),
  .c_addr_8_14(c_addr_8_14),
  .c_data_8_15(c_data_8_15),
  .c_addr_8_15(c_addr_8_15),
  .c_data_9_0(c_data_9_0),
  .c_addr_9_0(c_addr_9_0),
  .c_data_9_1(c_data_9_1),
  .c_addr_9_1(c_addr_9_1),
  .c_data_9_2(c_data_9_2),
  .c_addr_9_2(c_addr_9_2),
  .c_data_9_3(c_data_9_3),
  .c_addr_9_3(c_addr_9_3),
  .c_data_9_4(c_data_9_4),
  .c_addr_9_4(c_addr_9_4),
  .c_data_9_5(c_data_9_5),
  .c_addr_9_5(c_addr_9_5),
  .c_data_9_6(c_data_9_6),
  .c_addr_9_6(c_addr_9_6),
  .c_data_9_7(c_data_9_7),
  .c_addr_9_7(c_addr_9_7),
  .c_data_9_8(c_data_9_8),
  .c_addr_9_8(c_addr_9_8),
  .c_data_9_9(c_data_9_9),
  .c_addr_9_9(c_addr_9_9),
  .c_data_9_10(c_data_9_10),
  .c_addr_9_10(c_addr_9_10),
  .c_data_9_11(c_data_9_11),
  .c_addr_9_11(c_addr_9_11),
  .c_data_9_12(c_data_9_12),
  .c_addr_9_12(c_addr_9_12),
  .c_data_9_13(c_data_9_13),
  .c_addr_9_13(c_addr_9_13),
  .c_data_9_14(c_data_9_14),
  .c_addr_9_14(c_addr_9_14),
  .c_data_9_15(c_data_9_15),
  .c_addr_9_15(c_addr_9_15),
  .c_data_10_0(c_data_10_0),
  .c_addr_10_0(c_addr_10_0),
  .c_data_10_1(c_data_10_1),
  .c_addr_10_1(c_addr_10_1),
  .c_data_10_2(c_data_10_2),
  .c_addr_10_2(c_addr_10_2),
  .c_data_10_3(c_data_10_3),
  .c_addr_10_3(c_addr_10_3),
  .c_data_10_4(c_data_10_4),
  .c_addr_10_4(c_addr_10_4),
  .c_data_10_5(c_data_10_5),
  .c_addr_10_5(c_addr_10_5),
  .c_data_10_6(c_data_10_6),
  .c_addr_10_6(c_addr_10_6),
  .c_data_10_7(c_data_10_7),
  .c_addr_10_7(c_addr_10_7),
  .c_data_10_8(c_data_10_8),
  .c_addr_10_8(c_addr_10_8),
  .c_data_10_9(c_data_10_9),
  .c_addr_10_9(c_addr_10_9),
  .c_data_10_10(c_data_10_10),
  .c_addr_10_10(c_addr_10_10),
  .c_data_10_11(c_data_10_11),
  .c_addr_10_11(c_addr_10_11),
  .c_data_10_12(c_data_10_12),
  .c_addr_10_12(c_addr_10_12),
  .c_data_10_13(c_data_10_13),
  .c_addr_10_13(c_addr_10_13),
  .c_data_10_14(c_data_10_14),
  .c_addr_10_14(c_addr_10_14),
  .c_data_10_15(c_data_10_15),
  .c_addr_10_15(c_addr_10_15),
  .c_data_11_0(c_data_11_0),
  .c_addr_11_0(c_addr_11_0),
  .c_data_11_1(c_data_11_1),
  .c_addr_11_1(c_addr_11_1),
  .c_data_11_2(c_data_11_2),
  .c_addr_11_2(c_addr_11_2),
  .c_data_11_3(c_data_11_3),
  .c_addr_11_3(c_addr_11_3),
  .c_data_11_4(c_data_11_4),
  .c_addr_11_4(c_addr_11_4),
  .c_data_11_5(c_data_11_5),
  .c_addr_11_5(c_addr_11_5),
  .c_data_11_6(c_data_11_6),
  .c_addr_11_6(c_addr_11_6),
  .c_data_11_7(c_data_11_7),
  .c_addr_11_7(c_addr_11_7),
  .c_data_11_8(c_data_11_8),
  .c_addr_11_8(c_addr_11_8),
  .c_data_11_9(c_data_11_9),
  .c_addr_11_9(c_addr_11_9),
  .c_data_11_10(c_data_11_10),
  .c_addr_11_10(c_addr_11_10),
  .c_data_11_11(c_data_11_11),
  .c_addr_11_11(c_addr_11_11),
  .c_data_11_12(c_data_11_12),
  .c_addr_11_12(c_addr_11_12),
  .c_data_11_13(c_data_11_13),
  .c_addr_11_13(c_addr_11_13),
  .c_data_11_14(c_data_11_14),
  .c_addr_11_14(c_addr_11_14),
  .c_data_11_15(c_data_11_15),
  .c_addr_11_15(c_addr_11_15),
  .c_data_12_0(c_data_12_0),
  .c_addr_12_0(c_addr_12_0),
  .c_data_12_1(c_data_12_1),
  .c_addr_12_1(c_addr_12_1),
  .c_data_12_2(c_data_12_2),
  .c_addr_12_2(c_addr_12_2),
  .c_data_12_3(c_data_12_3),
  .c_addr_12_3(c_addr_12_3),
  .c_data_12_4(c_data_12_4),
  .c_addr_12_4(c_addr_12_4),
  .c_data_12_5(c_data_12_5),
  .c_addr_12_5(c_addr_12_5),
  .c_data_12_6(c_data_12_6),
  .c_addr_12_6(c_addr_12_6),
  .c_data_12_7(c_data_12_7),
  .c_addr_12_7(c_addr_12_7),
  .c_data_12_8(c_data_12_8),
  .c_addr_12_8(c_addr_12_8),
  .c_data_12_9(c_data_12_9),
  .c_addr_12_9(c_addr_12_9),
  .c_data_12_10(c_data_12_10),
  .c_addr_12_10(c_addr_12_10),
  .c_data_12_11(c_data_12_11),
  .c_addr_12_11(c_addr_12_11),
  .c_data_12_12(c_data_12_12),
  .c_addr_12_12(c_addr_12_12),
  .c_data_12_13(c_data_12_13),
  .c_addr_12_13(c_addr_12_13),
  .c_data_12_14(c_data_12_14),
  .c_addr_12_14(c_addr_12_14),
  .c_data_12_15(c_data_12_15),
  .c_addr_12_15(c_addr_12_15),
  .c_data_13_0(c_data_13_0),
  .c_addr_13_0(c_addr_13_0),
  .c_data_13_1(c_data_13_1),
  .c_addr_13_1(c_addr_13_1),
  .c_data_13_2(c_data_13_2),
  .c_addr_13_2(c_addr_13_2),
  .c_data_13_3(c_data_13_3),
  .c_addr_13_3(c_addr_13_3),
  .c_data_13_4(c_data_13_4),
  .c_addr_13_4(c_addr_13_4),
  .c_data_13_5(c_data_13_5),
  .c_addr_13_5(c_addr_13_5),
  .c_data_13_6(c_data_13_6),
  .c_addr_13_6(c_addr_13_6),
  .c_data_13_7(c_data_13_7),
  .c_addr_13_7(c_addr_13_7),
  .c_data_13_8(c_data_13_8),
  .c_addr_13_8(c_addr_13_8),
  .c_data_13_9(c_data_13_9),
  .c_addr_13_9(c_addr_13_9),
  .c_data_13_10(c_data_13_10),
  .c_addr_13_10(c_addr_13_10),
  .c_data_13_11(c_data_13_11),
  .c_addr_13_11(c_addr_13_11),
  .c_data_13_12(c_data_13_12),
  .c_addr_13_12(c_addr_13_12),
  .c_data_13_13(c_data_13_13),
  .c_addr_13_13(c_addr_13_13),
  .c_data_13_14(c_data_13_14),
  .c_addr_13_14(c_addr_13_14),
  .c_data_13_15(c_data_13_15),
  .c_addr_13_15(c_addr_13_15),
  .c_data_14_0(c_data_14_0),
  .c_addr_14_0(c_addr_14_0),
  .c_data_14_1(c_data_14_1),
  .c_addr_14_1(c_addr_14_1),
  .c_data_14_2(c_data_14_2),
  .c_addr_14_2(c_addr_14_2),
  .c_data_14_3(c_data_14_3),
  .c_addr_14_3(c_addr_14_3),
  .c_data_14_4(c_data_14_4),
  .c_addr_14_4(c_addr_14_4),
  .c_data_14_5(c_data_14_5),
  .c_addr_14_5(c_addr_14_5),
  .c_data_14_6(c_data_14_6),
  .c_addr_14_6(c_addr_14_6),
  .c_data_14_7(c_data_14_7),
  .c_addr_14_7(c_addr_14_7),
  .c_data_14_8(c_data_14_8),
  .c_addr_14_8(c_addr_14_8),
  .c_data_14_9(c_data_14_9),
  .c_addr_14_9(c_addr_14_9),
  .c_data_14_10(c_data_14_10),
  .c_addr_14_10(c_addr_14_10),
  .c_data_14_11(c_data_14_11),
  .c_addr_14_11(c_addr_14_11),
  .c_data_14_12(c_data_14_12),
  .c_addr_14_12(c_addr_14_12),
  .c_data_14_13(c_data_14_13),
  .c_addr_14_13(c_addr_14_13),
  .c_data_14_14(c_data_14_14),
  .c_addr_14_14(c_addr_14_14),
  .c_data_14_15(c_data_14_15),
  .c_addr_14_15(c_addr_14_15),
  .c_data_15_0(c_data_15_0),
  .c_addr_15_0(c_addr_15_0),
  .c_data_15_1(c_data_15_1),
  .c_addr_15_1(c_addr_15_1),
  .c_data_15_2(c_data_15_2),
  .c_addr_15_2(c_addr_15_2),
  .c_data_15_3(c_data_15_3),
  .c_addr_15_3(c_addr_15_3),
  .c_data_15_4(c_data_15_4),
  .c_addr_15_4(c_addr_15_4),
  .c_data_15_5(c_data_15_5),
  .c_addr_15_5(c_addr_15_5),
  .c_data_15_6(c_data_15_6),
  .c_addr_15_6(c_addr_15_6),
  .c_data_15_7(c_data_15_7),
  .c_addr_15_7(c_addr_15_7),
  .c_data_15_8(c_data_15_8),
  .c_addr_15_8(c_addr_15_8),
  .c_data_15_9(c_data_15_9),
  .c_addr_15_9(c_addr_15_9),
  .c_data_15_10(c_data_15_10),
  .c_addr_15_10(c_addr_15_10),
  .c_data_15_11(c_data_15_11),
  .c_addr_15_11(c_addr_15_11),
  .c_data_15_12(c_data_15_12),
  .c_addr_15_12(c_addr_15_12),
  .c_data_15_13(c_data_15_13),
  .c_addr_15_13(c_addr_15_13),
  .c_data_15_14(c_data_15_14),
  .c_addr_15_14(c_addr_15_14),
  .c_data_15_15(c_data_15_15),
  .c_addr_15_15(c_addr_15_15)

);
endmodule


/////////////////////////////////////////////////
// The 64x64 matmul definition
/////////////////////////////////////////////////

module matmul_64x64_systolic(
  clk,
  reset,
  start_mat_mul,
  done_mat_mul,
  a_data_0_0,
  a_addr_0_0,
  b_data_0_0,
  b_addr_0_0,
  a_data_1_0,
  a_addr_1_0,
  b_data_0_1,
  b_addr_0_1,
  a_data_2_0,
  a_addr_2_0,
  b_data_0_2,
  b_addr_0_2,
  a_data_3_0,
  a_addr_3_0,
  b_data_0_3,
  b_addr_0_3,
  a_data_4_0,
  a_addr_4_0,
  b_data_0_4,
  b_addr_0_4,
  a_data_5_0,
  a_addr_5_0,
  b_data_0_5,
  b_addr_0_5,
  a_data_6_0,
  a_addr_6_0,
  b_data_0_6,
  b_addr_0_6,
  a_data_7_0,
  a_addr_7_0,
  b_data_0_7,
  b_addr_0_7,
  a_data_8_0,
  a_addr_8_0,
  b_data_0_8,
  b_addr_0_8,
  a_data_9_0,
  a_addr_9_0,
  b_data_0_9,
  b_addr_0_9,
  a_data_10_0,
  a_addr_10_0,
  b_data_0_10,
  b_addr_0_10,
  a_data_11_0,
  a_addr_11_0,
  b_data_0_11,
  b_addr_0_11,
  a_data_12_0,
  a_addr_12_0,
  b_data_0_12,
  b_addr_0_12,
  a_data_13_0,
  a_addr_13_0,
  b_data_0_13,
  b_addr_0_13,
  a_data_14_0,
  a_addr_14_0,
  b_data_0_14,
  b_addr_0_14,
  a_data_15_0,
  a_addr_15_0,
  b_data_0_15,
  b_addr_0_15,

  c_data_0_0,
  c_addr_0_0,
  c_data_0_1,
  c_addr_0_1,
  c_data_0_2,
  c_addr_0_2,
  c_data_0_3,
  c_addr_0_3,
  c_data_0_4,
  c_addr_0_4,
  c_data_0_5,
  c_addr_0_5,
  c_data_0_6,
  c_addr_0_6,
  c_data_0_7,
  c_addr_0_7,
  c_data_0_8,
  c_addr_0_8,
  c_data_0_9,
  c_addr_0_9,
  c_data_0_10,
  c_addr_0_10,
  c_data_0_11,
  c_addr_0_11,
  c_data_0_12,
  c_addr_0_12,
  c_data_0_13,
  c_addr_0_13,
  c_data_0_14,
  c_addr_0_14,
  c_data_0_15,
  c_addr_0_15,
  c_data_1_0,
  c_addr_1_0,
  c_data_1_1,
  c_addr_1_1,
  c_data_1_2,
  c_addr_1_2,
  c_data_1_3,
  c_addr_1_3,
  c_data_1_4,
  c_addr_1_4,
  c_data_1_5,
  c_addr_1_5,
  c_data_1_6,
  c_addr_1_6,
  c_data_1_7,
  c_addr_1_7,
  c_data_1_8,
  c_addr_1_8,
  c_data_1_9,
  c_addr_1_9,
  c_data_1_10,
  c_addr_1_10,
  c_data_1_11,
  c_addr_1_11,
  c_data_1_12,
  c_addr_1_12,
  c_data_1_13,
  c_addr_1_13,
  c_data_1_14,
  c_addr_1_14,
  c_data_1_15,
  c_addr_1_15,
  c_data_2_0,
  c_addr_2_0,
  c_data_2_1,
  c_addr_2_1,
  c_data_2_2,
  c_addr_2_2,
  c_data_2_3,
  c_addr_2_3,
  c_data_2_4,
  c_addr_2_4,
  c_data_2_5,
  c_addr_2_5,
  c_data_2_6,
  c_addr_2_6,
  c_data_2_7,
  c_addr_2_7,
  c_data_2_8,
  c_addr_2_8,
  c_data_2_9,
  c_addr_2_9,
  c_data_2_10,
  c_addr_2_10,
  c_data_2_11,
  c_addr_2_11,
  c_data_2_12,
  c_addr_2_12,
  c_data_2_13,
  c_addr_2_13,
  c_data_2_14,
  c_addr_2_14,
  c_data_2_15,
  c_addr_2_15,
  c_data_3_0,
  c_addr_3_0,
  c_data_3_1,
  c_addr_3_1,
  c_data_3_2,
  c_addr_3_2,
  c_data_3_3,
  c_addr_3_3,
  c_data_3_4,
  c_addr_3_4,
  c_data_3_5,
  c_addr_3_5,
  c_data_3_6,
  c_addr_3_6,
  c_data_3_7,
  c_addr_3_7,
  c_data_3_8,
  c_addr_3_8,
  c_data_3_9,
  c_addr_3_9,
  c_data_3_10,
  c_addr_3_10,
  c_data_3_11,
  c_addr_3_11,
  c_data_3_12,
  c_addr_3_12,
  c_data_3_13,
  c_addr_3_13,
  c_data_3_14,
  c_addr_3_14,
  c_data_3_15,
  c_addr_3_15,
  c_data_4_0,
  c_addr_4_0,
  c_data_4_1,
  c_addr_4_1,
  c_data_4_2,
  c_addr_4_2,
  c_data_4_3,
  c_addr_4_3,
  c_data_4_4,
  c_addr_4_4,
  c_data_4_5,
  c_addr_4_5,
  c_data_4_6,
  c_addr_4_6,
  c_data_4_7,
  c_addr_4_7,
  c_data_4_8,
  c_addr_4_8,
  c_data_4_9,
  c_addr_4_9,
  c_data_4_10,
  c_addr_4_10,
  c_data_4_11,
  c_addr_4_11,
  c_data_4_12,
  c_addr_4_12,
  c_data_4_13,
  c_addr_4_13,
  c_data_4_14,
  c_addr_4_14,
  c_data_4_15,
  c_addr_4_15,
  c_data_5_0,
  c_addr_5_0,
  c_data_5_1,
  c_addr_5_1,
  c_data_5_2,
  c_addr_5_2,
  c_data_5_3,
  c_addr_5_3,
  c_data_5_4,
  c_addr_5_4,
  c_data_5_5,
  c_addr_5_5,
  c_data_5_6,
  c_addr_5_6,
  c_data_5_7,
  c_addr_5_7,
  c_data_5_8,
  c_addr_5_8,
  c_data_5_9,
  c_addr_5_9,
  c_data_5_10,
  c_addr_5_10,
  c_data_5_11,
  c_addr_5_11,
  c_data_5_12,
  c_addr_5_12,
  c_data_5_13,
  c_addr_5_13,
  c_data_5_14,
  c_addr_5_14,
  c_data_5_15,
  c_addr_5_15,
  c_data_6_0,
  c_addr_6_0,
  c_data_6_1,
  c_addr_6_1,
  c_data_6_2,
  c_addr_6_2,
  c_data_6_3,
  c_addr_6_3,
  c_data_6_4,
  c_addr_6_4,
  c_data_6_5,
  c_addr_6_5,
  c_data_6_6,
  c_addr_6_6,
  c_data_6_7,
  c_addr_6_7,
  c_data_6_8,
  c_addr_6_8,
  c_data_6_9,
  c_addr_6_9,
  c_data_6_10,
  c_addr_6_10,
  c_data_6_11,
  c_addr_6_11,
  c_data_6_12,
  c_addr_6_12,
  c_data_6_13,
  c_addr_6_13,
  c_data_6_14,
  c_addr_6_14,
  c_data_6_15,
  c_addr_6_15,
  c_data_7_0,
  c_addr_7_0,
  c_data_7_1,
  c_addr_7_1,
  c_data_7_2,
  c_addr_7_2,
  c_data_7_3,
  c_addr_7_3,
  c_data_7_4,
  c_addr_7_4,
  c_data_7_5,
  c_addr_7_5,
  c_data_7_6,
  c_addr_7_6,
  c_data_7_7,
  c_addr_7_7,
  c_data_7_8,
  c_addr_7_8,
  c_data_7_9,
  c_addr_7_9,
  c_data_7_10,
  c_addr_7_10,
  c_data_7_11,
  c_addr_7_11,
  c_data_7_12,
  c_addr_7_12,
  c_data_7_13,
  c_addr_7_13,
  c_data_7_14,
  c_addr_7_14,
  c_data_7_15,
  c_addr_7_15,
  c_data_8_0,
  c_addr_8_0,
  c_data_8_1,
  c_addr_8_1,
  c_data_8_2,
  c_addr_8_2,
  c_data_8_3,
  c_addr_8_3,
  c_data_8_4,
  c_addr_8_4,
  c_data_8_5,
  c_addr_8_5,
  c_data_8_6,
  c_addr_8_6,
  c_data_8_7,
  c_addr_8_7,
  c_data_8_8,
  c_addr_8_8,
  c_data_8_9,
  c_addr_8_9,
  c_data_8_10,
  c_addr_8_10,
  c_data_8_11,
  c_addr_8_11,
  c_data_8_12,
  c_addr_8_12,
  c_data_8_13,
  c_addr_8_13,
  c_data_8_14,
  c_addr_8_14,
  c_data_8_15,
  c_addr_8_15,
  c_data_9_0,
  c_addr_9_0,
  c_data_9_1,
  c_addr_9_1,
  c_data_9_2,
  c_addr_9_2,
  c_data_9_3,
  c_addr_9_3,
  c_data_9_4,
  c_addr_9_4,
  c_data_9_5,
  c_addr_9_5,
  c_data_9_6,
  c_addr_9_6,
  c_data_9_7,
  c_addr_9_7,
  c_data_9_8,
  c_addr_9_8,
  c_data_9_9,
  c_addr_9_9,
  c_data_9_10,
  c_addr_9_10,
  c_data_9_11,
  c_addr_9_11,
  c_data_9_12,
  c_addr_9_12,
  c_data_9_13,
  c_addr_9_13,
  c_data_9_14,
  c_addr_9_14,
  c_data_9_15,
  c_addr_9_15,
  c_data_10_0,
  c_addr_10_0,
  c_data_10_1,
  c_addr_10_1,
  c_data_10_2,
  c_addr_10_2,
  c_data_10_3,
  c_addr_10_3,
  c_data_10_4,
  c_addr_10_4,
  c_data_10_5,
  c_addr_10_5,
  c_data_10_6,
  c_addr_10_6,
  c_data_10_7,
  c_addr_10_7,
  c_data_10_8,
  c_addr_10_8,
  c_data_10_9,
  c_addr_10_9,
  c_data_10_10,
  c_addr_10_10,
  c_data_10_11,
  c_addr_10_11,
  c_data_10_12,
  c_addr_10_12,
  c_data_10_13,
  c_addr_10_13,
  c_data_10_14,
  c_addr_10_14,
  c_data_10_15,
  c_addr_10_15,
  c_data_11_0,
  c_addr_11_0,
  c_data_11_1,
  c_addr_11_1,
  c_data_11_2,
  c_addr_11_2,
  c_data_11_3,
  c_addr_11_3,
  c_data_11_4,
  c_addr_11_4,
  c_data_11_5,
  c_addr_11_5,
  c_data_11_6,
  c_addr_11_6,
  c_data_11_7,
  c_addr_11_7,
  c_data_11_8,
  c_addr_11_8,
  c_data_11_9,
  c_addr_11_9,
  c_data_11_10,
  c_addr_11_10,
  c_data_11_11,
  c_addr_11_11,
  c_data_11_12,
  c_addr_11_12,
  c_data_11_13,
  c_addr_11_13,
  c_data_11_14,
  c_addr_11_14,
  c_data_11_15,
  c_addr_11_15,
  c_data_12_0,
  c_addr_12_0,
  c_data_12_1,
  c_addr_12_1,
  c_data_12_2,
  c_addr_12_2,
  c_data_12_3,
  c_addr_12_3,
  c_data_12_4,
  c_addr_12_4,
  c_data_12_5,
  c_addr_12_5,
  c_data_12_6,
  c_addr_12_6,
  c_data_12_7,
  c_addr_12_7,
  c_data_12_8,
  c_addr_12_8,
  c_data_12_9,
  c_addr_12_9,
  c_data_12_10,
  c_addr_12_10,
  c_data_12_11,
  c_addr_12_11,
  c_data_12_12,
  c_addr_12_12,
  c_data_12_13,
  c_addr_12_13,
  c_data_12_14,
  c_addr_12_14,
  c_data_12_15,
  c_addr_12_15,
  c_data_13_0,
  c_addr_13_0,
  c_data_13_1,
  c_addr_13_1,
  c_data_13_2,
  c_addr_13_2,
  c_data_13_3,
  c_addr_13_3,
  c_data_13_4,
  c_addr_13_4,
  c_data_13_5,
  c_addr_13_5,
  c_data_13_6,
  c_addr_13_6,
  c_data_13_7,
  c_addr_13_7,
  c_data_13_8,
  c_addr_13_8,
  c_data_13_9,
  c_addr_13_9,
  c_data_13_10,
  c_addr_13_10,
  c_data_13_11,
  c_addr_13_11,
  c_data_13_12,
  c_addr_13_12,
  c_data_13_13,
  c_addr_13_13,
  c_data_13_14,
  c_addr_13_14,
  c_data_13_15,
  c_addr_13_15,
  c_data_14_0,
  c_addr_14_0,
  c_data_14_1,
  c_addr_14_1,
  c_data_14_2,
  c_addr_14_2,
  c_data_14_3,
  c_addr_14_3,
  c_data_14_4,
  c_addr_14_4,
  c_data_14_5,
  c_addr_14_5,
  c_data_14_6,
  c_addr_14_6,
  c_data_14_7,
  c_addr_14_7,
  c_data_14_8,
  c_addr_14_8,
  c_data_14_9,
  c_addr_14_9,
  c_data_14_10,
  c_addr_14_10,
  c_data_14_11,
  c_addr_14_11,
  c_data_14_12,
  c_addr_14_12,
  c_data_14_13,
  c_addr_14_13,
  c_data_14_14,
  c_addr_14_14,
  c_data_14_15,
  c_addr_14_15,
  c_data_15_0,
  c_addr_15_0,
  c_data_15_1,
  c_addr_15_1,
  c_data_15_2,
  c_addr_15_2,
  c_data_15_3,
  c_addr_15_3,
  c_data_15_4,
  c_addr_15_4,
  c_data_15_5,
  c_addr_15_5,
  c_data_15_6,
  c_addr_15_6,
  c_data_15_7,
  c_addr_15_7,
  c_data_15_8,
  c_addr_15_8,
  c_data_15_9,
  c_addr_15_9,
  c_data_15_10,
  c_addr_15_10,
  c_data_15_11,
  c_addr_15_11,
  c_data_15_12,
  c_addr_15_12,
  c_data_15_13,
  c_addr_15_13,
  c_data_15_14,
  c_addr_15_14,
  c_data_15_15,
  c_addr_15_15
);
  input clk;
  input reset;
  input start_mat_mul;
  output done_mat_mul;

  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_0;

  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_0;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_1;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_2;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_3;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_4;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_5;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_6;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_7;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_8;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_9;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_10;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_11;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_12;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_13;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_14;
  input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_15;

  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_0_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_1_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_2_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_3_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_4_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_5_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_6_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_7_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_8_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_9_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_10_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_11_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_12_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_13_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_14_15;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_0;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_1;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_2;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_3;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_4;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_5;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_6;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_7;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_8;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_9;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_10;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_11;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_12;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_13;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_14;
  output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] c_data_15_15;

  output [`AWIDTH-1:0] a_addr_0_0;
  output [`AWIDTH-1:0] a_addr_1_0;
  output [`AWIDTH-1:0] a_addr_2_0;
  output [`AWIDTH-1:0] a_addr_3_0;
  output [`AWIDTH-1:0] a_addr_4_0;
  output [`AWIDTH-1:0] a_addr_5_0;
  output [`AWIDTH-1:0] a_addr_6_0;
  output [`AWIDTH-1:0] a_addr_7_0;
  output [`AWIDTH-1:0] a_addr_8_0;
  output [`AWIDTH-1:0] a_addr_9_0;
  output [`AWIDTH-1:0] a_addr_10_0;
  output [`AWIDTH-1:0] a_addr_11_0;
  output [`AWIDTH-1:0] a_addr_12_0;
  output [`AWIDTH-1:0] a_addr_13_0;
  output [`AWIDTH-1:0] a_addr_14_0;
  output [`AWIDTH-1:0] a_addr_15_0;

  output [`AWIDTH-1:0] b_addr_0_0;
  output [`AWIDTH-1:0] b_addr_0_1;
  output [`AWIDTH-1:0] b_addr_0_2;
  output [`AWIDTH-1:0] b_addr_0_3;
  output [`AWIDTH-1:0] b_addr_0_4;
  output [`AWIDTH-1:0] b_addr_0_5;
  output [`AWIDTH-1:0] b_addr_0_6;
  output [`AWIDTH-1:0] b_addr_0_7;
  output [`AWIDTH-1:0] b_addr_0_8;
  output [`AWIDTH-1:0] b_addr_0_9;
  output [`AWIDTH-1:0] b_addr_0_10;
  output [`AWIDTH-1:0] b_addr_0_11;
  output [`AWIDTH-1:0] b_addr_0_12;
  output [`AWIDTH-1:0] b_addr_0_13;
  output [`AWIDTH-1:0] b_addr_0_14;
  output [`AWIDTH-1:0] b_addr_0_15;

  output [`AWIDTH-1:0] c_addr_0_0;
  output [`AWIDTH-1:0] c_addr_0_1;
  output [`AWIDTH-1:0] c_addr_0_2;
  output [`AWIDTH-1:0] c_addr_0_3;
  output [`AWIDTH-1:0] c_addr_0_4;
  output [`AWIDTH-1:0] c_addr_0_5;
  output [`AWIDTH-1:0] c_addr_0_6;
  output [`AWIDTH-1:0] c_addr_0_7;
  output [`AWIDTH-1:0] c_addr_0_8;
  output [`AWIDTH-1:0] c_addr_0_9;
  output [`AWIDTH-1:0] c_addr_0_10;
  output [`AWIDTH-1:0] c_addr_0_11;
  output [`AWIDTH-1:0] c_addr_0_12;
  output [`AWIDTH-1:0] c_addr_0_13;
  output [`AWIDTH-1:0] c_addr_0_14;
  output [`AWIDTH-1:0] c_addr_0_15;
  output [`AWIDTH-1:0] c_addr_1_0;
  output [`AWIDTH-1:0] c_addr_1_1;
  output [`AWIDTH-1:0] c_addr_1_2;
  output [`AWIDTH-1:0] c_addr_1_3;
  output [`AWIDTH-1:0] c_addr_1_4;
  output [`AWIDTH-1:0] c_addr_1_5;
  output [`AWIDTH-1:0] c_addr_1_6;
  output [`AWIDTH-1:0] c_addr_1_7;
  output [`AWIDTH-1:0] c_addr_1_8;
  output [`AWIDTH-1:0] c_addr_1_9;
  output [`AWIDTH-1:0] c_addr_1_10;
  output [`AWIDTH-1:0] c_addr_1_11;
  output [`AWIDTH-1:0] c_addr_1_12;
  output [`AWIDTH-1:0] c_addr_1_13;
  output [`AWIDTH-1:0] c_addr_1_14;
  output [`AWIDTH-1:0] c_addr_1_15;
  output [`AWIDTH-1:0] c_addr_2_0;
  output [`AWIDTH-1:0] c_addr_2_1;
  output [`AWIDTH-1:0] c_addr_2_2;
  output [`AWIDTH-1:0] c_addr_2_3;
  output [`AWIDTH-1:0] c_addr_2_4;
  output [`AWIDTH-1:0] c_addr_2_5;
  output [`AWIDTH-1:0] c_addr_2_6;
  output [`AWIDTH-1:0] c_addr_2_7;
  output [`AWIDTH-1:0] c_addr_2_8;
  output [`AWIDTH-1:0] c_addr_2_9;
  output [`AWIDTH-1:0] c_addr_2_10;
  output [`AWIDTH-1:0] c_addr_2_11;
  output [`AWIDTH-1:0] c_addr_2_12;
  output [`AWIDTH-1:0] c_addr_2_13;
  output [`AWIDTH-1:0] c_addr_2_14;
  output [`AWIDTH-1:0] c_addr_2_15;
  output [`AWIDTH-1:0] c_addr_3_0;
  output [`AWIDTH-1:0] c_addr_3_1;
  output [`AWIDTH-1:0] c_addr_3_2;
  output [`AWIDTH-1:0] c_addr_3_3;
  output [`AWIDTH-1:0] c_addr_3_4;
  output [`AWIDTH-1:0] c_addr_3_5;
  output [`AWIDTH-1:0] c_addr_3_6;
  output [`AWIDTH-1:0] c_addr_3_7;
  output [`AWIDTH-1:0] c_addr_3_8;
  output [`AWIDTH-1:0] c_addr_3_9;
  output [`AWIDTH-1:0] c_addr_3_10;
  output [`AWIDTH-1:0] c_addr_3_11;
  output [`AWIDTH-1:0] c_addr_3_12;
  output [`AWIDTH-1:0] c_addr_3_13;
  output [`AWIDTH-1:0] c_addr_3_14;
  output [`AWIDTH-1:0] c_addr_3_15;
  output [`AWIDTH-1:0] c_addr_4_0;
  output [`AWIDTH-1:0] c_addr_4_1;
  output [`AWIDTH-1:0] c_addr_4_2;
  output [`AWIDTH-1:0] c_addr_4_3;
  output [`AWIDTH-1:0] c_addr_4_4;
  output [`AWIDTH-1:0] c_addr_4_5;
  output [`AWIDTH-1:0] c_addr_4_6;
  output [`AWIDTH-1:0] c_addr_4_7;
  output [`AWIDTH-1:0] c_addr_4_8;
  output [`AWIDTH-1:0] c_addr_4_9;
  output [`AWIDTH-1:0] c_addr_4_10;
  output [`AWIDTH-1:0] c_addr_4_11;
  output [`AWIDTH-1:0] c_addr_4_12;
  output [`AWIDTH-1:0] c_addr_4_13;
  output [`AWIDTH-1:0] c_addr_4_14;
  output [`AWIDTH-1:0] c_addr_4_15;
  output [`AWIDTH-1:0] c_addr_5_0;
  output [`AWIDTH-1:0] c_addr_5_1;
  output [`AWIDTH-1:0] c_addr_5_2;
  output [`AWIDTH-1:0] c_addr_5_3;
  output [`AWIDTH-1:0] c_addr_5_4;
  output [`AWIDTH-1:0] c_addr_5_5;
  output [`AWIDTH-1:0] c_addr_5_6;
  output [`AWIDTH-1:0] c_addr_5_7;
  output [`AWIDTH-1:0] c_addr_5_8;
  output [`AWIDTH-1:0] c_addr_5_9;
  output [`AWIDTH-1:0] c_addr_5_10;
  output [`AWIDTH-1:0] c_addr_5_11;
  output [`AWIDTH-1:0] c_addr_5_12;
  output [`AWIDTH-1:0] c_addr_5_13;
  output [`AWIDTH-1:0] c_addr_5_14;
  output [`AWIDTH-1:0] c_addr_5_15;
  output [`AWIDTH-1:0] c_addr_6_0;
  output [`AWIDTH-1:0] c_addr_6_1;
  output [`AWIDTH-1:0] c_addr_6_2;
  output [`AWIDTH-1:0] c_addr_6_3;
  output [`AWIDTH-1:0] c_addr_6_4;
  output [`AWIDTH-1:0] c_addr_6_5;
  output [`AWIDTH-1:0] c_addr_6_6;
  output [`AWIDTH-1:0] c_addr_6_7;
  output [`AWIDTH-1:0] c_addr_6_8;
  output [`AWIDTH-1:0] c_addr_6_9;
  output [`AWIDTH-1:0] c_addr_6_10;
  output [`AWIDTH-1:0] c_addr_6_11;
  output [`AWIDTH-1:0] c_addr_6_12;
  output [`AWIDTH-1:0] c_addr_6_13;
  output [`AWIDTH-1:0] c_addr_6_14;
  output [`AWIDTH-1:0] c_addr_6_15;
  output [`AWIDTH-1:0] c_addr_7_0;
  output [`AWIDTH-1:0] c_addr_7_1;
  output [`AWIDTH-1:0] c_addr_7_2;
  output [`AWIDTH-1:0] c_addr_7_3;
  output [`AWIDTH-1:0] c_addr_7_4;
  output [`AWIDTH-1:0] c_addr_7_5;
  output [`AWIDTH-1:0] c_addr_7_6;
  output [`AWIDTH-1:0] c_addr_7_7;
  output [`AWIDTH-1:0] c_addr_7_8;
  output [`AWIDTH-1:0] c_addr_7_9;
  output [`AWIDTH-1:0] c_addr_7_10;
  output [`AWIDTH-1:0] c_addr_7_11;
  output [`AWIDTH-1:0] c_addr_7_12;
  output [`AWIDTH-1:0] c_addr_7_13;
  output [`AWIDTH-1:0] c_addr_7_14;
  output [`AWIDTH-1:0] c_addr_7_15;
  output [`AWIDTH-1:0] c_addr_8_0;
  output [`AWIDTH-1:0] c_addr_8_1;
  output [`AWIDTH-1:0] c_addr_8_2;
  output [`AWIDTH-1:0] c_addr_8_3;
  output [`AWIDTH-1:0] c_addr_8_4;
  output [`AWIDTH-1:0] c_addr_8_5;
  output [`AWIDTH-1:0] c_addr_8_6;
  output [`AWIDTH-1:0] c_addr_8_7;
  output [`AWIDTH-1:0] c_addr_8_8;
  output [`AWIDTH-1:0] c_addr_8_9;
  output [`AWIDTH-1:0] c_addr_8_10;
  output [`AWIDTH-1:0] c_addr_8_11;
  output [`AWIDTH-1:0] c_addr_8_12;
  output [`AWIDTH-1:0] c_addr_8_13;
  output [`AWIDTH-1:0] c_addr_8_14;
  output [`AWIDTH-1:0] c_addr_8_15;
  output [`AWIDTH-1:0] c_addr_9_0;
  output [`AWIDTH-1:0] c_addr_9_1;
  output [`AWIDTH-1:0] c_addr_9_2;
  output [`AWIDTH-1:0] c_addr_9_3;
  output [`AWIDTH-1:0] c_addr_9_4;
  output [`AWIDTH-1:0] c_addr_9_5;
  output [`AWIDTH-1:0] c_addr_9_6;
  output [`AWIDTH-1:0] c_addr_9_7;
  output [`AWIDTH-1:0] c_addr_9_8;
  output [`AWIDTH-1:0] c_addr_9_9;
  output [`AWIDTH-1:0] c_addr_9_10;
  output [`AWIDTH-1:0] c_addr_9_11;
  output [`AWIDTH-1:0] c_addr_9_12;
  output [`AWIDTH-1:0] c_addr_9_13;
  output [`AWIDTH-1:0] c_addr_9_14;
  output [`AWIDTH-1:0] c_addr_9_15;
  output [`AWIDTH-1:0] c_addr_10_0;
  output [`AWIDTH-1:0] c_addr_10_1;
  output [`AWIDTH-1:0] c_addr_10_2;
  output [`AWIDTH-1:0] c_addr_10_3;
  output [`AWIDTH-1:0] c_addr_10_4;
  output [`AWIDTH-1:0] c_addr_10_5;
  output [`AWIDTH-1:0] c_addr_10_6;
  output [`AWIDTH-1:0] c_addr_10_7;
  output [`AWIDTH-1:0] c_addr_10_8;
  output [`AWIDTH-1:0] c_addr_10_9;
  output [`AWIDTH-1:0] c_addr_10_10;
  output [`AWIDTH-1:0] c_addr_10_11;
  output [`AWIDTH-1:0] c_addr_10_12;
  output [`AWIDTH-1:0] c_addr_10_13;
  output [`AWIDTH-1:0] c_addr_10_14;
  output [`AWIDTH-1:0] c_addr_10_15;
  output [`AWIDTH-1:0] c_addr_11_0;
  output [`AWIDTH-1:0] c_addr_11_1;
  output [`AWIDTH-1:0] c_addr_11_2;
  output [`AWIDTH-1:0] c_addr_11_3;
  output [`AWIDTH-1:0] c_addr_11_4;
  output [`AWIDTH-1:0] c_addr_11_5;
  output [`AWIDTH-1:0] c_addr_11_6;
  output [`AWIDTH-1:0] c_addr_11_7;
  output [`AWIDTH-1:0] c_addr_11_8;
  output [`AWIDTH-1:0] c_addr_11_9;
  output [`AWIDTH-1:0] c_addr_11_10;
  output [`AWIDTH-1:0] c_addr_11_11;
  output [`AWIDTH-1:0] c_addr_11_12;
  output [`AWIDTH-1:0] c_addr_11_13;
  output [`AWIDTH-1:0] c_addr_11_14;
  output [`AWIDTH-1:0] c_addr_11_15;
  output [`AWIDTH-1:0] c_addr_12_0;
  output [`AWIDTH-1:0] c_addr_12_1;
  output [`AWIDTH-1:0] c_addr_12_2;
  output [`AWIDTH-1:0] c_addr_12_3;
  output [`AWIDTH-1:0] c_addr_12_4;
  output [`AWIDTH-1:0] c_addr_12_5;
  output [`AWIDTH-1:0] c_addr_12_6;
  output [`AWIDTH-1:0] c_addr_12_7;
  output [`AWIDTH-1:0] c_addr_12_8;
  output [`AWIDTH-1:0] c_addr_12_9;
  output [`AWIDTH-1:0] c_addr_12_10;
  output [`AWIDTH-1:0] c_addr_12_11;
  output [`AWIDTH-1:0] c_addr_12_12;
  output [`AWIDTH-1:0] c_addr_12_13;
  output [`AWIDTH-1:0] c_addr_12_14;
  output [`AWIDTH-1:0] c_addr_12_15;
  output [`AWIDTH-1:0] c_addr_13_0;
  output [`AWIDTH-1:0] c_addr_13_1;
  output [`AWIDTH-1:0] c_addr_13_2;
  output [`AWIDTH-1:0] c_addr_13_3;
  output [`AWIDTH-1:0] c_addr_13_4;
  output [`AWIDTH-1:0] c_addr_13_5;
  output [`AWIDTH-1:0] c_addr_13_6;
  output [`AWIDTH-1:0] c_addr_13_7;
  output [`AWIDTH-1:0] c_addr_13_8;
  output [`AWIDTH-1:0] c_addr_13_9;
  output [`AWIDTH-1:0] c_addr_13_10;
  output [`AWIDTH-1:0] c_addr_13_11;
  output [`AWIDTH-1:0] c_addr_13_12;
  output [`AWIDTH-1:0] c_addr_13_13;
  output [`AWIDTH-1:0] c_addr_13_14;
  output [`AWIDTH-1:0] c_addr_13_15;
  output [`AWIDTH-1:0] c_addr_14_0;
  output [`AWIDTH-1:0] c_addr_14_1;
  output [`AWIDTH-1:0] c_addr_14_2;
  output [`AWIDTH-1:0] c_addr_14_3;
  output [`AWIDTH-1:0] c_addr_14_4;
  output [`AWIDTH-1:0] c_addr_14_5;
  output [`AWIDTH-1:0] c_addr_14_6;
  output [`AWIDTH-1:0] c_addr_14_7;
  output [`AWIDTH-1:0] c_addr_14_8;
  output [`AWIDTH-1:0] c_addr_14_9;
  output [`AWIDTH-1:0] c_addr_14_10;
  output [`AWIDTH-1:0] c_addr_14_11;
  output [`AWIDTH-1:0] c_addr_14_12;
  output [`AWIDTH-1:0] c_addr_14_13;
  output [`AWIDTH-1:0] c_addr_14_14;
  output [`AWIDTH-1:0] c_addr_14_15;
  output [`AWIDTH-1:0] c_addr_15_0;
  output [`AWIDTH-1:0] c_addr_15_1;
  output [`AWIDTH-1:0] c_addr_15_2;
  output [`AWIDTH-1:0] c_addr_15_3;
  output [`AWIDTH-1:0] c_addr_15_4;
  output [`AWIDTH-1:0] c_addr_15_5;
  output [`AWIDTH-1:0] c_addr_15_6;
  output [`AWIDTH-1:0] c_addr_15_7;
  output [`AWIDTH-1:0] c_addr_15_8;
  output [`AWIDTH-1:0] c_addr_15_9;
  output [`AWIDTH-1:0] c_addr_15_10;
  output [`AWIDTH-1:0] c_addr_15_11;
  output [`AWIDTH-1:0] c_addr_15_12;
  output [`AWIDTH-1:0] c_addr_15_13;
  output [`AWIDTH-1:0] c_addr_15_14;
  output [`AWIDTH-1:0] c_addr_15_15;

  /////////////////////////////////////////////////
  // ORing all done signals
  /////////////////////////////////////////////////
  wire done_mat_mul_0_0;
  wire done_mat_mul_0_1;
  wire done_mat_mul_0_2;
  wire done_mat_mul_0_3;
  wire done_mat_mul_0_4;
  wire done_mat_mul_0_5;
  wire done_mat_mul_0_6;
  wire done_mat_mul_0_7;
  wire done_mat_mul_0_8;
  wire done_mat_mul_0_9;
  wire done_mat_mul_0_10;
  wire done_mat_mul_0_11;
  wire done_mat_mul_0_12;
  wire done_mat_mul_0_13;
  wire done_mat_mul_0_14;
  wire done_mat_mul_0_15;
  wire done_mat_mul_1_0;
  wire done_mat_mul_1_1;
  wire done_mat_mul_1_2;
  wire done_mat_mul_1_3;
  wire done_mat_mul_1_4;
  wire done_mat_mul_1_5;
  wire done_mat_mul_1_6;
  wire done_mat_mul_1_7;
  wire done_mat_mul_1_8;
  wire done_mat_mul_1_9;
  wire done_mat_mul_1_10;
  wire done_mat_mul_1_11;
  wire done_mat_mul_1_12;
  wire done_mat_mul_1_13;
  wire done_mat_mul_1_14;
  wire done_mat_mul_1_15;
  wire done_mat_mul_2_0;
  wire done_mat_mul_2_1;
  wire done_mat_mul_2_2;
  wire done_mat_mul_2_3;
  wire done_mat_mul_2_4;
  wire done_mat_mul_2_5;
  wire done_mat_mul_2_6;
  wire done_mat_mul_2_7;
  wire done_mat_mul_2_8;
  wire done_mat_mul_2_9;
  wire done_mat_mul_2_10;
  wire done_mat_mul_2_11;
  wire done_mat_mul_2_12;
  wire done_mat_mul_2_13;
  wire done_mat_mul_2_14;
  wire done_mat_mul_2_15;
  wire done_mat_mul_3_0;
  wire done_mat_mul_3_1;
  wire done_mat_mul_3_2;
  wire done_mat_mul_3_3;
  wire done_mat_mul_3_4;
  wire done_mat_mul_3_5;
  wire done_mat_mul_3_6;
  wire done_mat_mul_3_7;
  wire done_mat_mul_3_8;
  wire done_mat_mul_3_9;
  wire done_mat_mul_3_10;
  wire done_mat_mul_3_11;
  wire done_mat_mul_3_12;
  wire done_mat_mul_3_13;
  wire done_mat_mul_3_14;
  wire done_mat_mul_3_15;
  wire done_mat_mul_4_0;
  wire done_mat_mul_4_1;
  wire done_mat_mul_4_2;
  wire done_mat_mul_4_3;
  wire done_mat_mul_4_4;
  wire done_mat_mul_4_5;
  wire done_mat_mul_4_6;
  wire done_mat_mul_4_7;
  wire done_mat_mul_4_8;
  wire done_mat_mul_4_9;
  wire done_mat_mul_4_10;
  wire done_mat_mul_4_11;
  wire done_mat_mul_4_12;
  wire done_mat_mul_4_13;
  wire done_mat_mul_4_14;
  wire done_mat_mul_4_15;
  wire done_mat_mul_5_0;
  wire done_mat_mul_5_1;
  wire done_mat_mul_5_2;
  wire done_mat_mul_5_3;
  wire done_mat_mul_5_4;
  wire done_mat_mul_5_5;
  wire done_mat_mul_5_6;
  wire done_mat_mul_5_7;
  wire done_mat_mul_5_8;
  wire done_mat_mul_5_9;
  wire done_mat_mul_5_10;
  wire done_mat_mul_5_11;
  wire done_mat_mul_5_12;
  wire done_mat_mul_5_13;
  wire done_mat_mul_5_14;
  wire done_mat_mul_5_15;
  wire done_mat_mul_6_0;
  wire done_mat_mul_6_1;
  wire done_mat_mul_6_2;
  wire done_mat_mul_6_3;
  wire done_mat_mul_6_4;
  wire done_mat_mul_6_5;
  wire done_mat_mul_6_6;
  wire done_mat_mul_6_7;
  wire done_mat_mul_6_8;
  wire done_mat_mul_6_9;
  wire done_mat_mul_6_10;
  wire done_mat_mul_6_11;
  wire done_mat_mul_6_12;
  wire done_mat_mul_6_13;
  wire done_mat_mul_6_14;
  wire done_mat_mul_6_15;
  wire done_mat_mul_7_0;
  wire done_mat_mul_7_1;
  wire done_mat_mul_7_2;
  wire done_mat_mul_7_3;
  wire done_mat_mul_7_4;
  wire done_mat_mul_7_5;
  wire done_mat_mul_7_6;
  wire done_mat_mul_7_7;
  wire done_mat_mul_7_8;
  wire done_mat_mul_7_9;
  wire done_mat_mul_7_10;
  wire done_mat_mul_7_11;
  wire done_mat_mul_7_12;
  wire done_mat_mul_7_13;
  wire done_mat_mul_7_14;
  wire done_mat_mul_7_15;
  wire done_mat_mul_8_0;
  wire done_mat_mul_8_1;
  wire done_mat_mul_8_2;
  wire done_mat_mul_8_3;
  wire done_mat_mul_8_4;
  wire done_mat_mul_8_5;
  wire done_mat_mul_8_6;
  wire done_mat_mul_8_7;
  wire done_mat_mul_8_8;
  wire done_mat_mul_8_9;
  wire done_mat_mul_8_10;
  wire done_mat_mul_8_11;
  wire done_mat_mul_8_12;
  wire done_mat_mul_8_13;
  wire done_mat_mul_8_14;
  wire done_mat_mul_8_15;
  wire done_mat_mul_9_0;
  wire done_mat_mul_9_1;
  wire done_mat_mul_9_2;
  wire done_mat_mul_9_3;
  wire done_mat_mul_9_4;
  wire done_mat_mul_9_5;
  wire done_mat_mul_9_6;
  wire done_mat_mul_9_7;
  wire done_mat_mul_9_8;
  wire done_mat_mul_9_9;
  wire done_mat_mul_9_10;
  wire done_mat_mul_9_11;
  wire done_mat_mul_9_12;
  wire done_mat_mul_9_13;
  wire done_mat_mul_9_14;
  wire done_mat_mul_9_15;
  wire done_mat_mul_10_0;
  wire done_mat_mul_10_1;
  wire done_mat_mul_10_2;
  wire done_mat_mul_10_3;
  wire done_mat_mul_10_4;
  wire done_mat_mul_10_5;
  wire done_mat_mul_10_6;
  wire done_mat_mul_10_7;
  wire done_mat_mul_10_8;
  wire done_mat_mul_10_9;
  wire done_mat_mul_10_10;
  wire done_mat_mul_10_11;
  wire done_mat_mul_10_12;
  wire done_mat_mul_10_13;
  wire done_mat_mul_10_14;
  wire done_mat_mul_10_15;
  wire done_mat_mul_11_0;
  wire done_mat_mul_11_1;
  wire done_mat_mul_11_2;
  wire done_mat_mul_11_3;
  wire done_mat_mul_11_4;
  wire done_mat_mul_11_5;
  wire done_mat_mul_11_6;
  wire done_mat_mul_11_7;
  wire done_mat_mul_11_8;
  wire done_mat_mul_11_9;
  wire done_mat_mul_11_10;
  wire done_mat_mul_11_11;
  wire done_mat_mul_11_12;
  wire done_mat_mul_11_13;
  wire done_mat_mul_11_14;
  wire done_mat_mul_11_15;
  wire done_mat_mul_12_0;
  wire done_mat_mul_12_1;
  wire done_mat_mul_12_2;
  wire done_mat_mul_12_3;
  wire done_mat_mul_12_4;
  wire done_mat_mul_12_5;
  wire done_mat_mul_12_6;
  wire done_mat_mul_12_7;
  wire done_mat_mul_12_8;
  wire done_mat_mul_12_9;
  wire done_mat_mul_12_10;
  wire done_mat_mul_12_11;
  wire done_mat_mul_12_12;
  wire done_mat_mul_12_13;
  wire done_mat_mul_12_14;
  wire done_mat_mul_12_15;
  wire done_mat_mul_13_0;
  wire done_mat_mul_13_1;
  wire done_mat_mul_13_2;
  wire done_mat_mul_13_3;
  wire done_mat_mul_13_4;
  wire done_mat_mul_13_5;
  wire done_mat_mul_13_6;
  wire done_mat_mul_13_7;
  wire done_mat_mul_13_8;
  wire done_mat_mul_13_9;
  wire done_mat_mul_13_10;
  wire done_mat_mul_13_11;
  wire done_mat_mul_13_12;
  wire done_mat_mul_13_13;
  wire done_mat_mul_13_14;
  wire done_mat_mul_13_15;
  wire done_mat_mul_14_0;
  wire done_mat_mul_14_1;
  wire done_mat_mul_14_2;
  wire done_mat_mul_14_3;
  wire done_mat_mul_14_4;
  wire done_mat_mul_14_5;
  wire done_mat_mul_14_6;
  wire done_mat_mul_14_7;
  wire done_mat_mul_14_8;
  wire done_mat_mul_14_9;
  wire done_mat_mul_14_10;
  wire done_mat_mul_14_11;
  wire done_mat_mul_14_12;
  wire done_mat_mul_14_13;
  wire done_mat_mul_14_14;
  wire done_mat_mul_14_15;
  wire done_mat_mul_15_0;
  wire done_mat_mul_15_1;
  wire done_mat_mul_15_2;
  wire done_mat_mul_15_3;
  wire done_mat_mul_15_4;
  wire done_mat_mul_15_5;
  wire done_mat_mul_15_6;
  wire done_mat_mul_15_7;
  wire done_mat_mul_15_8;
  wire done_mat_mul_15_9;
  wire done_mat_mul_15_10;
  wire done_mat_mul_15_11;
  wire done_mat_mul_15_12;
  wire done_mat_mul_15_13;
  wire done_mat_mul_15_14;
  wire done_mat_mul_15_15;

  assign done_mat_mul =   done_mat_mul_0_0 &&
  done_mat_mul_0_1 &&
  done_mat_mul_0_2 &&
  done_mat_mul_0_3 &&
  done_mat_mul_0_4 &&
  done_mat_mul_0_5 &&
  done_mat_mul_0_6 &&
  done_mat_mul_0_7 &&
  done_mat_mul_0_8 &&
  done_mat_mul_0_9 &&
  done_mat_mul_0_10 &&
  done_mat_mul_0_11 &&
  done_mat_mul_0_12 &&
  done_mat_mul_0_13 &&
  done_mat_mul_0_14 &&
  done_mat_mul_0_15 &&
  done_mat_mul_1_0 &&
  done_mat_mul_1_1 &&
  done_mat_mul_1_2 &&
  done_mat_mul_1_3 &&
  done_mat_mul_1_4 &&
  done_mat_mul_1_5 &&
  done_mat_mul_1_6 &&
  done_mat_mul_1_7 &&
  done_mat_mul_1_8 &&
  done_mat_mul_1_9 &&
  done_mat_mul_1_10 &&
  done_mat_mul_1_11 &&
  done_mat_mul_1_12 &&
  done_mat_mul_1_13 &&
  done_mat_mul_1_14 &&
  done_mat_mul_1_15 &&
  done_mat_mul_2_0 &&
  done_mat_mul_2_1 &&
  done_mat_mul_2_2 &&
  done_mat_mul_2_3 &&
  done_mat_mul_2_4 &&
  done_mat_mul_2_5 &&
  done_mat_mul_2_6 &&
  done_mat_mul_2_7 &&
  done_mat_mul_2_8 &&
  done_mat_mul_2_9 &&
  done_mat_mul_2_10 &&
  done_mat_mul_2_11 &&
  done_mat_mul_2_12 &&
  done_mat_mul_2_13 &&
  done_mat_mul_2_14 &&
  done_mat_mul_2_15 &&
  done_mat_mul_3_0 &&
  done_mat_mul_3_1 &&
  done_mat_mul_3_2 &&
  done_mat_mul_3_3 &&
  done_mat_mul_3_4 &&
  done_mat_mul_3_5 &&
  done_mat_mul_3_6 &&
  done_mat_mul_3_7 &&
  done_mat_mul_3_8 &&
  done_mat_mul_3_9 &&
  done_mat_mul_3_10 &&
  done_mat_mul_3_11 &&
  done_mat_mul_3_12 &&
  done_mat_mul_3_13 &&
  done_mat_mul_3_14 &&
  done_mat_mul_3_15 &&
  done_mat_mul_4_0 &&
  done_mat_mul_4_1 &&
  done_mat_mul_4_2 &&
  done_mat_mul_4_3 &&
  done_mat_mul_4_4 &&
  done_mat_mul_4_5 &&
  done_mat_mul_4_6 &&
  done_mat_mul_4_7 &&
  done_mat_mul_4_8 &&
  done_mat_mul_4_9 &&
  done_mat_mul_4_10 &&
  done_mat_mul_4_11 &&
  done_mat_mul_4_12 &&
  done_mat_mul_4_13 &&
  done_mat_mul_4_14 &&
  done_mat_mul_4_15 &&
  done_mat_mul_5_0 &&
  done_mat_mul_5_1 &&
  done_mat_mul_5_2 &&
  done_mat_mul_5_3 &&
  done_mat_mul_5_4 &&
  done_mat_mul_5_5 &&
  done_mat_mul_5_6 &&
  done_mat_mul_5_7 &&
  done_mat_mul_5_8 &&
  done_mat_mul_5_9 &&
  done_mat_mul_5_10 &&
  done_mat_mul_5_11 &&
  done_mat_mul_5_12 &&
  done_mat_mul_5_13 &&
  done_mat_mul_5_14 &&
  done_mat_mul_5_15 &&
  done_mat_mul_6_0 &&
  done_mat_mul_6_1 &&
  done_mat_mul_6_2 &&
  done_mat_mul_6_3 &&
  done_mat_mul_6_4 &&
  done_mat_mul_6_5 &&
  done_mat_mul_6_6 &&
  done_mat_mul_6_7 &&
  done_mat_mul_6_8 &&
  done_mat_mul_6_9 &&
  done_mat_mul_6_10 &&
  done_mat_mul_6_11 &&
  done_mat_mul_6_12 &&
  done_mat_mul_6_13 &&
  done_mat_mul_6_14 &&
  done_mat_mul_6_15 &&
  done_mat_mul_7_0 &&
  done_mat_mul_7_1 &&
  done_mat_mul_7_2 &&
  done_mat_mul_7_3 &&
  done_mat_mul_7_4 &&
  done_mat_mul_7_5 &&
  done_mat_mul_7_6 &&
  done_mat_mul_7_7 &&
  done_mat_mul_7_8 &&
  done_mat_mul_7_9 &&
  done_mat_mul_7_10 &&
  done_mat_mul_7_11 &&
  done_mat_mul_7_12 &&
  done_mat_mul_7_13 &&
  done_mat_mul_7_14 &&
  done_mat_mul_7_15 &&
  done_mat_mul_8_0 &&
  done_mat_mul_8_1 &&
  done_mat_mul_8_2 &&
  done_mat_mul_8_3 &&
  done_mat_mul_8_4 &&
  done_mat_mul_8_5 &&
  done_mat_mul_8_6 &&
  done_mat_mul_8_7 &&
  done_mat_mul_8_8 &&
  done_mat_mul_8_9 &&
  done_mat_mul_8_10 &&
  done_mat_mul_8_11 &&
  done_mat_mul_8_12 &&
  done_mat_mul_8_13 &&
  done_mat_mul_8_14 &&
  done_mat_mul_8_15 &&
  done_mat_mul_9_0 &&
  done_mat_mul_9_1 &&
  done_mat_mul_9_2 &&
  done_mat_mul_9_3 &&
  done_mat_mul_9_4 &&
  done_mat_mul_9_5 &&
  done_mat_mul_9_6 &&
  done_mat_mul_9_7 &&
  done_mat_mul_9_8 &&
  done_mat_mul_9_9 &&
  done_mat_mul_9_10 &&
  done_mat_mul_9_11 &&
  done_mat_mul_9_12 &&
  done_mat_mul_9_13 &&
  done_mat_mul_9_14 &&
  done_mat_mul_9_15 &&
  done_mat_mul_10_0 &&
  done_mat_mul_10_1 &&
  done_mat_mul_10_2 &&
  done_mat_mul_10_3 &&
  done_mat_mul_10_4 &&
  done_mat_mul_10_5 &&
  done_mat_mul_10_6 &&
  done_mat_mul_10_7 &&
  done_mat_mul_10_8 &&
  done_mat_mul_10_9 &&
  done_mat_mul_10_10 &&
  done_mat_mul_10_11 &&
  done_mat_mul_10_12 &&
  done_mat_mul_10_13 &&
  done_mat_mul_10_14 &&
  done_mat_mul_10_15 &&
  done_mat_mul_11_0 &&
  done_mat_mul_11_1 &&
  done_mat_mul_11_2 &&
  done_mat_mul_11_3 &&
  done_mat_mul_11_4 &&
  done_mat_mul_11_5 &&
  done_mat_mul_11_6 &&
  done_mat_mul_11_7 &&
  done_mat_mul_11_8 &&
  done_mat_mul_11_9 &&
  done_mat_mul_11_10 &&
  done_mat_mul_11_11 &&
  done_mat_mul_11_12 &&
  done_mat_mul_11_13 &&
  done_mat_mul_11_14 &&
  done_mat_mul_11_15 &&
  done_mat_mul_12_0 &&
  done_mat_mul_12_1 &&
  done_mat_mul_12_2 &&
  done_mat_mul_12_3 &&
  done_mat_mul_12_4 &&
  done_mat_mul_12_5 &&
  done_mat_mul_12_6 &&
  done_mat_mul_12_7 &&
  done_mat_mul_12_8 &&
  done_mat_mul_12_9 &&
  done_mat_mul_12_10 &&
  done_mat_mul_12_11 &&
  done_mat_mul_12_12 &&
  done_mat_mul_12_13 &&
  done_mat_mul_12_14 &&
  done_mat_mul_12_15 &&
  done_mat_mul_13_0 &&
  done_mat_mul_13_1 &&
  done_mat_mul_13_2 &&
  done_mat_mul_13_3 &&
  done_mat_mul_13_4 &&
  done_mat_mul_13_5 &&
  done_mat_mul_13_6 &&
  done_mat_mul_13_7 &&
  done_mat_mul_13_8 &&
  done_mat_mul_13_9 &&
  done_mat_mul_13_10 &&
  done_mat_mul_13_11 &&
  done_mat_mul_13_12 &&
  done_mat_mul_13_13 &&
  done_mat_mul_13_14 &&
  done_mat_mul_13_15 &&
  done_mat_mul_14_0 &&
  done_mat_mul_14_1 &&
  done_mat_mul_14_2 &&
  done_mat_mul_14_3 &&
  done_mat_mul_14_4 &&
  done_mat_mul_14_5 &&
  done_mat_mul_14_6 &&
  done_mat_mul_14_7 &&
  done_mat_mul_14_8 &&
  done_mat_mul_14_9 &&
  done_mat_mul_14_10 &&
  done_mat_mul_14_11 &&
  done_mat_mul_14_12 &&
  done_mat_mul_14_13 &&
  done_mat_mul_14_14 &&
  done_mat_mul_14_15 &&
  done_mat_mul_15_0 &&
  done_mat_mul_15_1 &&
  done_mat_mul_15_2 &&
  done_mat_mul_15_3 &&
  done_mat_mul_15_4 &&
  done_mat_mul_15_5 &&
  done_mat_mul_15_6 &&
  done_mat_mul_15_7 &&
  done_mat_mul_15_8 &&
  done_mat_mul_15_9 &&
  done_mat_mul_15_10 &&
  done_mat_mul_15_11 &&
  done_mat_mul_15_12 &&
  done_mat_mul_15_13 &&
  done_mat_mul_15_14 &&
  done_mat_mul_15_15;

  /////////////////////////////////////////////////
  // Matmul 0_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_0_to_0_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_0_to_1_0;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_0_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_0),
  .a_data(a_data_0_0),
  .b_data(b_data_0_0),
  .a_data_in(a_data_in_0_0_NC),
  .b_data_in(b_data_in_0_0_NC),
  .c_data(c_data_0_0),
  .a_data_out(a_data_0_0_to_0_1),
  .b_data_out(b_data_0_0_to_1_0),
  .a_addr(a_addr_0_0),
  .b_addr(b_addr_0_0),
  .c_addr(c_addr_0_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 0_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_1_to_0_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_1_to_1_1;
  wire [`AWIDTH-1:0] a_addr_0_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_1),
  .a_data(a_data_0_1_NC),
  .b_data(b_data_0_1),
  .a_data_in(a_data_0_0_to_0_1),
  .b_data_in(b_data_in_0_1_NC),
  .c_data(c_data_0_1),
  .a_data_out(a_data_0_1_to_0_2),
  .b_data_out(b_data_0_1_to_1_1),
  .a_addr(a_addr_0_1_NC),
  .b_addr(b_addr_0_1),
  .c_addr(c_addr_0_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 0_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_2_to_0_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_2_to_1_2;
  wire [`AWIDTH-1:0] a_addr_0_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_2),
  .a_data(a_data_0_2_NC),
  .b_data(b_data_0_2),
  .a_data_in(a_data_0_1_to_0_2),
  .b_data_in(b_data_in_0_2_NC),
  .c_data(c_data_0_2),
  .a_data_out(a_data_0_2_to_0_3),
  .b_data_out(b_data_0_2_to_1_2),
  .a_addr(a_addr_0_2_NC),
  .b_addr(b_addr_0_2),
  .c_addr(c_addr_0_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 0_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_3_to_0_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_3_to_1_3;
  wire [`AWIDTH-1:0] a_addr_0_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_3),
  .a_data(a_data_0_3_NC),
  .b_data(b_data_0_3),
  .a_data_in(a_data_0_2_to_0_3),
  .b_data_in(b_data_in_0_3_NC),
  .c_data(c_data_0_3),
  .a_data_out(a_data_0_3_to_0_4),
  .b_data_out(b_data_0_3_to_1_3),
  .a_addr(a_addr_0_3_NC),
  .b_addr(b_addr_0_3),
  .c_addr(c_addr_0_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 0_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_4_to_0_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_4_to_1_4;
  wire [`AWIDTH-1:0] a_addr_0_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_4),
  .a_data(a_data_0_4_NC),
  .b_data(b_data_0_4),
  .a_data_in(a_data_0_3_to_0_4),
  .b_data_in(b_data_in_0_4_NC),
  .c_data(c_data_0_4),
  .a_data_out(a_data_0_4_to_0_5),
  .b_data_out(b_data_0_4_to_1_4),
  .a_addr(a_addr_0_4_NC),
  .b_addr(b_addr_0_4),
  .c_addr(c_addr_0_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 0_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_5_to_0_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_5_to_1_5;
  wire [`AWIDTH-1:0] a_addr_0_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_5),
  .a_data(a_data_0_5_NC),
  .b_data(b_data_0_5),
  .a_data_in(a_data_0_4_to_0_5),
  .b_data_in(b_data_in_0_5_NC),
  .c_data(c_data_0_5),
  .a_data_out(a_data_0_5_to_0_6),
  .b_data_out(b_data_0_5_to_1_5),
  .a_addr(a_addr_0_5_NC),
  .b_addr(b_addr_0_5),
  .c_addr(c_addr_0_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 0_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_6_to_0_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_6_to_1_6;
  wire [`AWIDTH-1:0] a_addr_0_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_6),
  .a_data(a_data_0_6_NC),
  .b_data(b_data_0_6),
  .a_data_in(a_data_0_5_to_0_6),
  .b_data_in(b_data_in_0_6_NC),
  .c_data(c_data_0_6),
  .a_data_out(a_data_0_6_to_0_7),
  .b_data_out(b_data_0_6_to_1_6),
  .a_addr(a_addr_0_6_NC),
  .b_addr(b_addr_0_6),
  .c_addr(c_addr_0_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 0_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_7_to_0_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_7_to_1_7;
  wire [`AWIDTH-1:0] a_addr_0_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_7),
  .a_data(a_data_0_7_NC),
  .b_data(b_data_0_7),
  .a_data_in(a_data_0_6_to_0_7),
  .b_data_in(b_data_in_0_7_NC),
  .c_data(c_data_0_7),
  .a_data_out(a_data_0_7_to_0_8),
  .b_data_out(b_data_0_7_to_1_7),
  .a_addr(a_addr_0_7_NC),
  .b_addr(b_addr_0_7),
  .c_addr(c_addr_0_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 0_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_8_to_0_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_8_to_1_8;
  wire [`AWIDTH-1:0] a_addr_0_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_8),
  .a_data(a_data_0_8_NC),
  .b_data(b_data_0_8),
  .a_data_in(a_data_0_7_to_0_8),
  .b_data_in(b_data_in_0_8_NC),
  .c_data(c_data_0_8),
  .a_data_out(a_data_0_8_to_0_9),
  .b_data_out(b_data_0_8_to_1_8),
  .a_addr(a_addr_0_8_NC),
  .b_addr(b_addr_0_8),
  .c_addr(c_addr_0_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 0_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_9_to_0_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_9_to_1_9;
  wire [`AWIDTH-1:0] a_addr_0_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_9),
  .a_data(a_data_0_9_NC),
  .b_data(b_data_0_9),
  .a_data_in(a_data_0_8_to_0_9),
  .b_data_in(b_data_in_0_9_NC),
  .c_data(c_data_0_9),
  .a_data_out(a_data_0_9_to_0_10),
  .b_data_out(b_data_0_9_to_1_9),
  .a_addr(a_addr_0_9_NC),
  .b_addr(b_addr_0_9),
  .c_addr(c_addr_0_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 0_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_10_to_0_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_10_to_1_10;
  wire [`AWIDTH-1:0] a_addr_0_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_10),
  .a_data(a_data_0_10_NC),
  .b_data(b_data_0_10),
  .a_data_in(a_data_0_9_to_0_10),
  .b_data_in(b_data_in_0_10_NC),
  .c_data(c_data_0_10),
  .a_data_out(a_data_0_10_to_0_11),
  .b_data_out(b_data_0_10_to_1_10),
  .a_addr(a_addr_0_10_NC),
  .b_addr(b_addr_0_10),
  .c_addr(c_addr_0_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 0_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_11_to_0_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_11_to_1_11;
  wire [`AWIDTH-1:0] a_addr_0_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_11),
  .a_data(a_data_0_11_NC),
  .b_data(b_data_0_11),
  .a_data_in(a_data_0_10_to_0_11),
  .b_data_in(b_data_in_0_11_NC),
  .c_data(c_data_0_11),
  .a_data_out(a_data_0_11_to_0_12),
  .b_data_out(b_data_0_11_to_1_11),
  .a_addr(a_addr_0_11_NC),
  .b_addr(b_addr_0_11),
  .c_addr(c_addr_0_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 0_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_12_to_0_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_12_to_1_12;
  wire [`AWIDTH-1:0] a_addr_0_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_12),
  .a_data(a_data_0_12_NC),
  .b_data(b_data_0_12),
  .a_data_in(a_data_0_11_to_0_12),
  .b_data_in(b_data_in_0_12_NC),
  .c_data(c_data_0_12),
  .a_data_out(a_data_0_12_to_0_13),
  .b_data_out(b_data_0_12_to_1_12),
  .a_addr(a_addr_0_12_NC),
  .b_addr(b_addr_0_12),
  .c_addr(c_addr_0_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 0_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_13_to_0_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_13_to_1_13;
  wire [`AWIDTH-1:0] a_addr_0_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_13),
  .a_data(a_data_0_13_NC),
  .b_data(b_data_0_13),
  .a_data_in(a_data_0_12_to_0_13),
  .b_data_in(b_data_in_0_13_NC),
  .c_data(c_data_0_13),
  .a_data_out(a_data_0_13_to_0_14),
  .b_data_out(b_data_0_13_to_1_13),
  .a_addr(a_addr_0_13_NC),
  .b_addr(b_addr_0_13),
  .c_addr(c_addr_0_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 0_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_14_to_0_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_14_to_1_14;
  wire [`AWIDTH-1:0] a_addr_0_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_14),
  .a_data(a_data_0_14_NC),
  .b_data(b_data_0_14),
  .a_data_in(a_data_0_13_to_0_14),
  .b_data_in(b_data_in_0_14_NC),
  .c_data(c_data_0_14),
  .a_data_out(a_data_0_14_to_0_15),
  .b_data_out(b_data_0_14_to_1_14),
  .a_addr(a_addr_0_14_NC),
  .b_addr(b_addr_0_14),
  .c_addr(c_addr_0_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 0_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_15_to_0_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_0_15_to_1_15;
  wire [`AWIDTH-1:0] a_addr_0_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_0_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in_0_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_0_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_0_15),
  .a_data(a_data_0_15_NC),
  .b_data(b_data_0_15),
  .a_data_in(a_data_0_14_to_0_15),
  .b_data_in(b_data_in_0_15_NC),
  .c_data(c_data_0_15),
  .a_data_out(a_data_0_15_to_0_16),
  .b_data_out(b_data_0_15_to_1_15),
  .a_addr(a_addr_0_15_NC),
  .b_addr(b_addr_0_15),
  .c_addr(c_addr_0_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd0),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 1_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_0_to_1_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_0_to_2_0;
  wire [`AWIDTH-1:0] b_addr_1_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_1_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_0),
  .a_data(a_data_1_0),
  .b_data(b_data_1_0_NC),
  .a_data_in(a_data_in_1_0_NC),
  .b_data_in(b_data_0_0_to_1_0),
  .c_data(c_data_1_0),
  .a_data_out(a_data_1_0_to_1_1),
  .b_data_out(b_data_1_0_to_2_0),
  .a_addr(a_addr_1_0),
  .b_addr(b_addr_1_0_NC),
  .c_addr(c_addr_1_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 1_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_1_to_1_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_1_to_2_1;
  wire [`AWIDTH-1:0] a_addr_1_1_NC;
  wire [`AWIDTH-1:0] b_addr_1_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_1),
  .a_data(a_data_1_1_NC),
  .b_data(b_data_1_1_NC),
  .a_data_in(a_data_1_0_to_1_1),
  .b_data_in(b_data_0_1_to_1_1),
  .c_data(c_data_1_1),
  .a_data_out(a_data_1_1_to_1_2),
  .b_data_out(b_data_1_1_to_2_1),
  .a_addr(a_addr_1_1_NC),
  .b_addr(b_addr_1_1_NC),
  .c_addr(c_addr_1_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 1_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_2_to_1_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_2_to_2_2;
  wire [`AWIDTH-1:0] a_addr_1_2_NC;
  wire [`AWIDTH-1:0] b_addr_1_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_2),
  .a_data(a_data_1_2_NC),
  .b_data(b_data_1_2_NC),
  .a_data_in(a_data_1_1_to_1_2),
  .b_data_in(b_data_0_2_to_1_2),
  .c_data(c_data_1_2),
  .a_data_out(a_data_1_2_to_1_3),
  .b_data_out(b_data_1_2_to_2_2),
  .a_addr(a_addr_1_2_NC),
  .b_addr(b_addr_1_2_NC),
  .c_addr(c_addr_1_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 1_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_3_to_1_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_3_to_2_3;
  wire [`AWIDTH-1:0] a_addr_1_3_NC;
  wire [`AWIDTH-1:0] b_addr_1_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_3),
  .a_data(a_data_1_3_NC),
  .b_data(b_data_1_3_NC),
  .a_data_in(a_data_1_2_to_1_3),
  .b_data_in(b_data_0_3_to_1_3),
  .c_data(c_data_1_3),
  .a_data_out(a_data_1_3_to_1_4),
  .b_data_out(b_data_1_3_to_2_3),
  .a_addr(a_addr_1_3_NC),
  .b_addr(b_addr_1_3_NC),
  .c_addr(c_addr_1_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 1_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_4_to_1_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_4_to_2_4;
  wire [`AWIDTH-1:0] a_addr_1_4_NC;
  wire [`AWIDTH-1:0] b_addr_1_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_4),
  .a_data(a_data_1_4_NC),
  .b_data(b_data_1_4_NC),
  .a_data_in(a_data_1_3_to_1_4),
  .b_data_in(b_data_0_4_to_1_4),
  .c_data(c_data_1_4),
  .a_data_out(a_data_1_4_to_1_5),
  .b_data_out(b_data_1_4_to_2_4),
  .a_addr(a_addr_1_4_NC),
  .b_addr(b_addr_1_4_NC),
  .c_addr(c_addr_1_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 1_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_5_to_1_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_5_to_2_5;
  wire [`AWIDTH-1:0] a_addr_1_5_NC;
  wire [`AWIDTH-1:0] b_addr_1_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_5),
  .a_data(a_data_1_5_NC),
  .b_data(b_data_1_5_NC),
  .a_data_in(a_data_1_4_to_1_5),
  .b_data_in(b_data_0_5_to_1_5),
  .c_data(c_data_1_5),
  .a_data_out(a_data_1_5_to_1_6),
  .b_data_out(b_data_1_5_to_2_5),
  .a_addr(a_addr_1_5_NC),
  .b_addr(b_addr_1_5_NC),
  .c_addr(c_addr_1_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 1_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_6_to_1_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_6_to_2_6;
  wire [`AWIDTH-1:0] a_addr_1_6_NC;
  wire [`AWIDTH-1:0] b_addr_1_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_6),
  .a_data(a_data_1_6_NC),
  .b_data(b_data_1_6_NC),
  .a_data_in(a_data_1_5_to_1_6),
  .b_data_in(b_data_0_6_to_1_6),
  .c_data(c_data_1_6),
  .a_data_out(a_data_1_6_to_1_7),
  .b_data_out(b_data_1_6_to_2_6),
  .a_addr(a_addr_1_6_NC),
  .b_addr(b_addr_1_6_NC),
  .c_addr(c_addr_1_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 1_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_7_to_1_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_7_to_2_7;
  wire [`AWIDTH-1:0] a_addr_1_7_NC;
  wire [`AWIDTH-1:0] b_addr_1_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_7),
  .a_data(a_data_1_7_NC),
  .b_data(b_data_1_7_NC),
  .a_data_in(a_data_1_6_to_1_7),
  .b_data_in(b_data_0_7_to_1_7),
  .c_data(c_data_1_7),
  .a_data_out(a_data_1_7_to_1_8),
  .b_data_out(b_data_1_7_to_2_7),
  .a_addr(a_addr_1_7_NC),
  .b_addr(b_addr_1_7_NC),
  .c_addr(c_addr_1_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 1_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_8_to_1_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_8_to_2_8;
  wire [`AWIDTH-1:0] a_addr_1_8_NC;
  wire [`AWIDTH-1:0] b_addr_1_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_8),
  .a_data(a_data_1_8_NC),
  .b_data(b_data_1_8_NC),
  .a_data_in(a_data_1_7_to_1_8),
  .b_data_in(b_data_0_8_to_1_8),
  .c_data(c_data_1_8),
  .a_data_out(a_data_1_8_to_1_9),
  .b_data_out(b_data_1_8_to_2_8),
  .a_addr(a_addr_1_8_NC),
  .b_addr(b_addr_1_8_NC),
  .c_addr(c_addr_1_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 1_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_9_to_1_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_9_to_2_9;
  wire [`AWIDTH-1:0] a_addr_1_9_NC;
  wire [`AWIDTH-1:0] b_addr_1_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_9),
  .a_data(a_data_1_9_NC),
  .b_data(b_data_1_9_NC),
  .a_data_in(a_data_1_8_to_1_9),
  .b_data_in(b_data_0_9_to_1_9),
  .c_data(c_data_1_9),
  .a_data_out(a_data_1_9_to_1_10),
  .b_data_out(b_data_1_9_to_2_9),
  .a_addr(a_addr_1_9_NC),
  .b_addr(b_addr_1_9_NC),
  .c_addr(c_addr_1_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 1_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_10_to_1_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_10_to_2_10;
  wire [`AWIDTH-1:0] a_addr_1_10_NC;
  wire [`AWIDTH-1:0] b_addr_1_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_10),
  .a_data(a_data_1_10_NC),
  .b_data(b_data_1_10_NC),
  .a_data_in(a_data_1_9_to_1_10),
  .b_data_in(b_data_0_10_to_1_10),
  .c_data(c_data_1_10),
  .a_data_out(a_data_1_10_to_1_11),
  .b_data_out(b_data_1_10_to_2_10),
  .a_addr(a_addr_1_10_NC),
  .b_addr(b_addr_1_10_NC),
  .c_addr(c_addr_1_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 1_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_11_to_1_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_11_to_2_11;
  wire [`AWIDTH-1:0] a_addr_1_11_NC;
  wire [`AWIDTH-1:0] b_addr_1_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_11),
  .a_data(a_data_1_11_NC),
  .b_data(b_data_1_11_NC),
  .a_data_in(a_data_1_10_to_1_11),
  .b_data_in(b_data_0_11_to_1_11),
  .c_data(c_data_1_11),
  .a_data_out(a_data_1_11_to_1_12),
  .b_data_out(b_data_1_11_to_2_11),
  .a_addr(a_addr_1_11_NC),
  .b_addr(b_addr_1_11_NC),
  .c_addr(c_addr_1_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 1_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_12_to_1_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_12_to_2_12;
  wire [`AWIDTH-1:0] a_addr_1_12_NC;
  wire [`AWIDTH-1:0] b_addr_1_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_12),
  .a_data(a_data_1_12_NC),
  .b_data(b_data_1_12_NC),
  .a_data_in(a_data_1_11_to_1_12),
  .b_data_in(b_data_0_12_to_1_12),
  .c_data(c_data_1_12),
  .a_data_out(a_data_1_12_to_1_13),
  .b_data_out(b_data_1_12_to_2_12),
  .a_addr(a_addr_1_12_NC),
  .b_addr(b_addr_1_12_NC),
  .c_addr(c_addr_1_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 1_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_13_to_1_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_13_to_2_13;
  wire [`AWIDTH-1:0] a_addr_1_13_NC;
  wire [`AWIDTH-1:0] b_addr_1_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_13),
  .a_data(a_data_1_13_NC),
  .b_data(b_data_1_13_NC),
  .a_data_in(a_data_1_12_to_1_13),
  .b_data_in(b_data_0_13_to_1_13),
  .c_data(c_data_1_13),
  .a_data_out(a_data_1_13_to_1_14),
  .b_data_out(b_data_1_13_to_2_13),
  .a_addr(a_addr_1_13_NC),
  .b_addr(b_addr_1_13_NC),
  .c_addr(c_addr_1_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 1_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_14_to_1_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_14_to_2_14;
  wire [`AWIDTH-1:0] a_addr_1_14_NC;
  wire [`AWIDTH-1:0] b_addr_1_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_14),
  .a_data(a_data_1_14_NC),
  .b_data(b_data_1_14_NC),
  .a_data_in(a_data_1_13_to_1_14),
  .b_data_in(b_data_0_14_to_1_14),
  .c_data(c_data_1_14),
  .a_data_out(a_data_1_14_to_1_15),
  .b_data_out(b_data_1_14_to_2_14),
  .a_addr(a_addr_1_14_NC),
  .b_addr(b_addr_1_14_NC),
  .c_addr(c_addr_1_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 1_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_15_to_1_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_15_to_2_15;
  wire [`AWIDTH-1:0] a_addr_1_15_NC;
  wire [`AWIDTH-1:0] b_addr_1_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_1_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_1_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_1_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_1_15),
  .a_data(a_data_1_15_NC),
  .b_data(b_data_1_15_NC),
  .a_data_in(a_data_1_14_to_1_15),
  .b_data_in(b_data_0_15_to_1_15),
  .c_data(c_data_1_15),
  .a_data_out(a_data_1_15_to_1_16),
  .b_data_out(b_data_1_15_to_2_15),
  .a_addr(a_addr_1_15_NC),
  .b_addr(b_addr_1_15_NC),
  .c_addr(c_addr_1_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd1),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 2_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_0_to_2_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_0_to_3_0;
  wire [`AWIDTH-1:0] b_addr_2_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_2_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_0),
  .a_data(a_data_2_0),
  .b_data(b_data_2_0_NC),
  .a_data_in(a_data_in_2_0_NC),
  .b_data_in(b_data_1_0_to_2_0),
  .c_data(c_data_2_0),
  .a_data_out(a_data_2_0_to_2_1),
  .b_data_out(b_data_2_0_to_3_0),
  .a_addr(a_addr_2_0),
  .b_addr(b_addr_2_0_NC),
  .c_addr(c_addr_2_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 2_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_1_to_2_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_1_to_3_1;
  wire [`AWIDTH-1:0] a_addr_2_1_NC;
  wire [`AWIDTH-1:0] b_addr_2_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_1),
  .a_data(a_data_2_1_NC),
  .b_data(b_data_2_1_NC),
  .a_data_in(a_data_2_0_to_2_1),
  .b_data_in(b_data_1_1_to_2_1),
  .c_data(c_data_2_1),
  .a_data_out(a_data_2_1_to_2_2),
  .b_data_out(b_data_2_1_to_3_1),
  .a_addr(a_addr_2_1_NC),
  .b_addr(b_addr_2_1_NC),
  .c_addr(c_addr_2_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 2_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_2_to_2_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_2_to_3_2;
  wire [`AWIDTH-1:0] a_addr_2_2_NC;
  wire [`AWIDTH-1:0] b_addr_2_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_2),
  .a_data(a_data_2_2_NC),
  .b_data(b_data_2_2_NC),
  .a_data_in(a_data_2_1_to_2_2),
  .b_data_in(b_data_1_2_to_2_2),
  .c_data(c_data_2_2),
  .a_data_out(a_data_2_2_to_2_3),
  .b_data_out(b_data_2_2_to_3_2),
  .a_addr(a_addr_2_2_NC),
  .b_addr(b_addr_2_2_NC),
  .c_addr(c_addr_2_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 2_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_3_to_2_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_3_to_3_3;
  wire [`AWIDTH-1:0] a_addr_2_3_NC;
  wire [`AWIDTH-1:0] b_addr_2_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_3),
  .a_data(a_data_2_3_NC),
  .b_data(b_data_2_3_NC),
  .a_data_in(a_data_2_2_to_2_3),
  .b_data_in(b_data_1_3_to_2_3),
  .c_data(c_data_2_3),
  .a_data_out(a_data_2_3_to_2_4),
  .b_data_out(b_data_2_3_to_3_3),
  .a_addr(a_addr_2_3_NC),
  .b_addr(b_addr_2_3_NC),
  .c_addr(c_addr_2_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 2_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_4_to_2_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_4_to_3_4;
  wire [`AWIDTH-1:0] a_addr_2_4_NC;
  wire [`AWIDTH-1:0] b_addr_2_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_4),
  .a_data(a_data_2_4_NC),
  .b_data(b_data_2_4_NC),
  .a_data_in(a_data_2_3_to_2_4),
  .b_data_in(b_data_1_4_to_2_4),
  .c_data(c_data_2_4),
  .a_data_out(a_data_2_4_to_2_5),
  .b_data_out(b_data_2_4_to_3_4),
  .a_addr(a_addr_2_4_NC),
  .b_addr(b_addr_2_4_NC),
  .c_addr(c_addr_2_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 2_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_5_to_2_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_5_to_3_5;
  wire [`AWIDTH-1:0] a_addr_2_5_NC;
  wire [`AWIDTH-1:0] b_addr_2_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_5),
  .a_data(a_data_2_5_NC),
  .b_data(b_data_2_5_NC),
  .a_data_in(a_data_2_4_to_2_5),
  .b_data_in(b_data_1_5_to_2_5),
  .c_data(c_data_2_5),
  .a_data_out(a_data_2_5_to_2_6),
  .b_data_out(b_data_2_5_to_3_5),
  .a_addr(a_addr_2_5_NC),
  .b_addr(b_addr_2_5_NC),
  .c_addr(c_addr_2_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 2_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_6_to_2_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_6_to_3_6;
  wire [`AWIDTH-1:0] a_addr_2_6_NC;
  wire [`AWIDTH-1:0] b_addr_2_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_6),
  .a_data(a_data_2_6_NC),
  .b_data(b_data_2_6_NC),
  .a_data_in(a_data_2_5_to_2_6),
  .b_data_in(b_data_1_6_to_2_6),
  .c_data(c_data_2_6),
  .a_data_out(a_data_2_6_to_2_7),
  .b_data_out(b_data_2_6_to_3_6),
  .a_addr(a_addr_2_6_NC),
  .b_addr(b_addr_2_6_NC),
  .c_addr(c_addr_2_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 2_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_7_to_2_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_7_to_3_7;
  wire [`AWIDTH-1:0] a_addr_2_7_NC;
  wire [`AWIDTH-1:0] b_addr_2_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_7),
  .a_data(a_data_2_7_NC),
  .b_data(b_data_2_7_NC),
  .a_data_in(a_data_2_6_to_2_7),
  .b_data_in(b_data_1_7_to_2_7),
  .c_data(c_data_2_7),
  .a_data_out(a_data_2_7_to_2_8),
  .b_data_out(b_data_2_7_to_3_7),
  .a_addr(a_addr_2_7_NC),
  .b_addr(b_addr_2_7_NC),
  .c_addr(c_addr_2_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 2_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_8_to_2_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_8_to_3_8;
  wire [`AWIDTH-1:0] a_addr_2_8_NC;
  wire [`AWIDTH-1:0] b_addr_2_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_8),
  .a_data(a_data_2_8_NC),
  .b_data(b_data_2_8_NC),
  .a_data_in(a_data_2_7_to_2_8),
  .b_data_in(b_data_1_8_to_2_8),
  .c_data(c_data_2_8),
  .a_data_out(a_data_2_8_to_2_9),
  .b_data_out(b_data_2_8_to_3_8),
  .a_addr(a_addr_2_8_NC),
  .b_addr(b_addr_2_8_NC),
  .c_addr(c_addr_2_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 2_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_9_to_2_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_9_to_3_9;
  wire [`AWIDTH-1:0] a_addr_2_9_NC;
  wire [`AWIDTH-1:0] b_addr_2_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_9),
  .a_data(a_data_2_9_NC),
  .b_data(b_data_2_9_NC),
  .a_data_in(a_data_2_8_to_2_9),
  .b_data_in(b_data_1_9_to_2_9),
  .c_data(c_data_2_9),
  .a_data_out(a_data_2_9_to_2_10),
  .b_data_out(b_data_2_9_to_3_9),
  .a_addr(a_addr_2_9_NC),
  .b_addr(b_addr_2_9_NC),
  .c_addr(c_addr_2_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 2_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_10_to_2_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_10_to_3_10;
  wire [`AWIDTH-1:0] a_addr_2_10_NC;
  wire [`AWIDTH-1:0] b_addr_2_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_10),
  .a_data(a_data_2_10_NC),
  .b_data(b_data_2_10_NC),
  .a_data_in(a_data_2_9_to_2_10),
  .b_data_in(b_data_1_10_to_2_10),
  .c_data(c_data_2_10),
  .a_data_out(a_data_2_10_to_2_11),
  .b_data_out(b_data_2_10_to_3_10),
  .a_addr(a_addr_2_10_NC),
  .b_addr(b_addr_2_10_NC),
  .c_addr(c_addr_2_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 2_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_11_to_2_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_11_to_3_11;
  wire [`AWIDTH-1:0] a_addr_2_11_NC;
  wire [`AWIDTH-1:0] b_addr_2_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_11),
  .a_data(a_data_2_11_NC),
  .b_data(b_data_2_11_NC),
  .a_data_in(a_data_2_10_to_2_11),
  .b_data_in(b_data_1_11_to_2_11),
  .c_data(c_data_2_11),
  .a_data_out(a_data_2_11_to_2_12),
  .b_data_out(b_data_2_11_to_3_11),
  .a_addr(a_addr_2_11_NC),
  .b_addr(b_addr_2_11_NC),
  .c_addr(c_addr_2_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 2_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_12_to_2_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_12_to_3_12;
  wire [`AWIDTH-1:0] a_addr_2_12_NC;
  wire [`AWIDTH-1:0] b_addr_2_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_12),
  .a_data(a_data_2_12_NC),
  .b_data(b_data_2_12_NC),
  .a_data_in(a_data_2_11_to_2_12),
  .b_data_in(b_data_1_12_to_2_12),
  .c_data(c_data_2_12),
  .a_data_out(a_data_2_12_to_2_13),
  .b_data_out(b_data_2_12_to_3_12),
  .a_addr(a_addr_2_12_NC),
  .b_addr(b_addr_2_12_NC),
  .c_addr(c_addr_2_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 2_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_13_to_2_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_13_to_3_13;
  wire [`AWIDTH-1:0] a_addr_2_13_NC;
  wire [`AWIDTH-1:0] b_addr_2_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_13),
  .a_data(a_data_2_13_NC),
  .b_data(b_data_2_13_NC),
  .a_data_in(a_data_2_12_to_2_13),
  .b_data_in(b_data_1_13_to_2_13),
  .c_data(c_data_2_13),
  .a_data_out(a_data_2_13_to_2_14),
  .b_data_out(b_data_2_13_to_3_13),
  .a_addr(a_addr_2_13_NC),
  .b_addr(b_addr_2_13_NC),
  .c_addr(c_addr_2_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 2_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_14_to_2_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_14_to_3_14;
  wire [`AWIDTH-1:0] a_addr_2_14_NC;
  wire [`AWIDTH-1:0] b_addr_2_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_14),
  .a_data(a_data_2_14_NC),
  .b_data(b_data_2_14_NC),
  .a_data_in(a_data_2_13_to_2_14),
  .b_data_in(b_data_1_14_to_2_14),
  .c_data(c_data_2_14),
  .a_data_out(a_data_2_14_to_2_15),
  .b_data_out(b_data_2_14_to_3_14),
  .a_addr(a_addr_2_14_NC),
  .b_addr(b_addr_2_14_NC),
  .c_addr(c_addr_2_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 2_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_15_to_2_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_15_to_3_15;
  wire [`AWIDTH-1:0] a_addr_2_15_NC;
  wire [`AWIDTH-1:0] b_addr_2_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_2_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_2_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_2_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_2_15),
  .a_data(a_data_2_15_NC),
  .b_data(b_data_2_15_NC),
  .a_data_in(a_data_2_14_to_2_15),
  .b_data_in(b_data_1_15_to_2_15),
  .c_data(c_data_2_15),
  .a_data_out(a_data_2_15_to_2_16),
  .b_data_out(b_data_2_15_to_3_15),
  .a_addr(a_addr_2_15_NC),
  .b_addr(b_addr_2_15_NC),
  .c_addr(c_addr_2_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd2),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 3_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_0_to_3_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_0_to_4_0;
  wire [`AWIDTH-1:0] b_addr_3_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_3_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_0),
  .a_data(a_data_3_0),
  .b_data(b_data_3_0_NC),
  .a_data_in(a_data_in_3_0_NC),
  .b_data_in(b_data_2_0_to_3_0),
  .c_data(c_data_3_0),
  .a_data_out(a_data_3_0_to_3_1),
  .b_data_out(b_data_3_0_to_4_0),
  .a_addr(a_addr_3_0),
  .b_addr(b_addr_3_0_NC),
  .c_addr(c_addr_3_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 3_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_1_to_3_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_1_to_4_1;
  wire [`AWIDTH-1:0] a_addr_3_1_NC;
  wire [`AWIDTH-1:0] b_addr_3_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_1),
  .a_data(a_data_3_1_NC),
  .b_data(b_data_3_1_NC),
  .a_data_in(a_data_3_0_to_3_1),
  .b_data_in(b_data_2_1_to_3_1),
  .c_data(c_data_3_1),
  .a_data_out(a_data_3_1_to_3_2),
  .b_data_out(b_data_3_1_to_4_1),
  .a_addr(a_addr_3_1_NC),
  .b_addr(b_addr_3_1_NC),
  .c_addr(c_addr_3_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 3_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_2_to_3_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_2_to_4_2;
  wire [`AWIDTH-1:0] a_addr_3_2_NC;
  wire [`AWIDTH-1:0] b_addr_3_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_2),
  .a_data(a_data_3_2_NC),
  .b_data(b_data_3_2_NC),
  .a_data_in(a_data_3_1_to_3_2),
  .b_data_in(b_data_2_2_to_3_2),
  .c_data(c_data_3_2),
  .a_data_out(a_data_3_2_to_3_3),
  .b_data_out(b_data_3_2_to_4_2),
  .a_addr(a_addr_3_2_NC),
  .b_addr(b_addr_3_2_NC),
  .c_addr(c_addr_3_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 3_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_3_to_3_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_3_to_4_3;
  wire [`AWIDTH-1:0] a_addr_3_3_NC;
  wire [`AWIDTH-1:0] b_addr_3_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_3),
  .a_data(a_data_3_3_NC),
  .b_data(b_data_3_3_NC),
  .a_data_in(a_data_3_2_to_3_3),
  .b_data_in(b_data_2_3_to_3_3),
  .c_data(c_data_3_3),
  .a_data_out(a_data_3_3_to_3_4),
  .b_data_out(b_data_3_3_to_4_3),
  .a_addr(a_addr_3_3_NC),
  .b_addr(b_addr_3_3_NC),
  .c_addr(c_addr_3_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 3_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_4_to_3_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_4_to_4_4;
  wire [`AWIDTH-1:0] a_addr_3_4_NC;
  wire [`AWIDTH-1:0] b_addr_3_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_4),
  .a_data(a_data_3_4_NC),
  .b_data(b_data_3_4_NC),
  .a_data_in(a_data_3_3_to_3_4),
  .b_data_in(b_data_2_4_to_3_4),
  .c_data(c_data_3_4),
  .a_data_out(a_data_3_4_to_3_5),
  .b_data_out(b_data_3_4_to_4_4),
  .a_addr(a_addr_3_4_NC),
  .b_addr(b_addr_3_4_NC),
  .c_addr(c_addr_3_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 3_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_5_to_3_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_5_to_4_5;
  wire [`AWIDTH-1:0] a_addr_3_5_NC;
  wire [`AWIDTH-1:0] b_addr_3_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_5),
  .a_data(a_data_3_5_NC),
  .b_data(b_data_3_5_NC),
  .a_data_in(a_data_3_4_to_3_5),
  .b_data_in(b_data_2_5_to_3_5),
  .c_data(c_data_3_5),
  .a_data_out(a_data_3_5_to_3_6),
  .b_data_out(b_data_3_5_to_4_5),
  .a_addr(a_addr_3_5_NC),
  .b_addr(b_addr_3_5_NC),
  .c_addr(c_addr_3_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 3_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_6_to_3_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_6_to_4_6;
  wire [`AWIDTH-1:0] a_addr_3_6_NC;
  wire [`AWIDTH-1:0] b_addr_3_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_6),
  .a_data(a_data_3_6_NC),
  .b_data(b_data_3_6_NC),
  .a_data_in(a_data_3_5_to_3_6),
  .b_data_in(b_data_2_6_to_3_6),
  .c_data(c_data_3_6),
  .a_data_out(a_data_3_6_to_3_7),
  .b_data_out(b_data_3_6_to_4_6),
  .a_addr(a_addr_3_6_NC),
  .b_addr(b_addr_3_6_NC),
  .c_addr(c_addr_3_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 3_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_7_to_3_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_7_to_4_7;
  wire [`AWIDTH-1:0] a_addr_3_7_NC;
  wire [`AWIDTH-1:0] b_addr_3_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_7),
  .a_data(a_data_3_7_NC),
  .b_data(b_data_3_7_NC),
  .a_data_in(a_data_3_6_to_3_7),
  .b_data_in(b_data_2_7_to_3_7),
  .c_data(c_data_3_7),
  .a_data_out(a_data_3_7_to_3_8),
  .b_data_out(b_data_3_7_to_4_7),
  .a_addr(a_addr_3_7_NC),
  .b_addr(b_addr_3_7_NC),
  .c_addr(c_addr_3_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 3_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_8_to_3_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_8_to_4_8;
  wire [`AWIDTH-1:0] a_addr_3_8_NC;
  wire [`AWIDTH-1:0] b_addr_3_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_8),
  .a_data(a_data_3_8_NC),
  .b_data(b_data_3_8_NC),
  .a_data_in(a_data_3_7_to_3_8),
  .b_data_in(b_data_2_8_to_3_8),
  .c_data(c_data_3_8),
  .a_data_out(a_data_3_8_to_3_9),
  .b_data_out(b_data_3_8_to_4_8),
  .a_addr(a_addr_3_8_NC),
  .b_addr(b_addr_3_8_NC),
  .c_addr(c_addr_3_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 3_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_9_to_3_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_9_to_4_9;
  wire [`AWIDTH-1:0] a_addr_3_9_NC;
  wire [`AWIDTH-1:0] b_addr_3_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_9),
  .a_data(a_data_3_9_NC),
  .b_data(b_data_3_9_NC),
  .a_data_in(a_data_3_8_to_3_9),
  .b_data_in(b_data_2_9_to_3_9),
  .c_data(c_data_3_9),
  .a_data_out(a_data_3_9_to_3_10),
  .b_data_out(b_data_3_9_to_4_9),
  .a_addr(a_addr_3_9_NC),
  .b_addr(b_addr_3_9_NC),
  .c_addr(c_addr_3_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 3_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_10_to_3_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_10_to_4_10;
  wire [`AWIDTH-1:0] a_addr_3_10_NC;
  wire [`AWIDTH-1:0] b_addr_3_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_10),
  .a_data(a_data_3_10_NC),
  .b_data(b_data_3_10_NC),
  .a_data_in(a_data_3_9_to_3_10),
  .b_data_in(b_data_2_10_to_3_10),
  .c_data(c_data_3_10),
  .a_data_out(a_data_3_10_to_3_11),
  .b_data_out(b_data_3_10_to_4_10),
  .a_addr(a_addr_3_10_NC),
  .b_addr(b_addr_3_10_NC),
  .c_addr(c_addr_3_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 3_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_11_to_3_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_11_to_4_11;
  wire [`AWIDTH-1:0] a_addr_3_11_NC;
  wire [`AWIDTH-1:0] b_addr_3_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_11),
  .a_data(a_data_3_11_NC),
  .b_data(b_data_3_11_NC),
  .a_data_in(a_data_3_10_to_3_11),
  .b_data_in(b_data_2_11_to_3_11),
  .c_data(c_data_3_11),
  .a_data_out(a_data_3_11_to_3_12),
  .b_data_out(b_data_3_11_to_4_11),
  .a_addr(a_addr_3_11_NC),
  .b_addr(b_addr_3_11_NC),
  .c_addr(c_addr_3_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 3_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_12_to_3_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_12_to_4_12;
  wire [`AWIDTH-1:0] a_addr_3_12_NC;
  wire [`AWIDTH-1:0] b_addr_3_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_12),
  .a_data(a_data_3_12_NC),
  .b_data(b_data_3_12_NC),
  .a_data_in(a_data_3_11_to_3_12),
  .b_data_in(b_data_2_12_to_3_12),
  .c_data(c_data_3_12),
  .a_data_out(a_data_3_12_to_3_13),
  .b_data_out(b_data_3_12_to_4_12),
  .a_addr(a_addr_3_12_NC),
  .b_addr(b_addr_3_12_NC),
  .c_addr(c_addr_3_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 3_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_13_to_3_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_13_to_4_13;
  wire [`AWIDTH-1:0] a_addr_3_13_NC;
  wire [`AWIDTH-1:0] b_addr_3_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_13),
  .a_data(a_data_3_13_NC),
  .b_data(b_data_3_13_NC),
  .a_data_in(a_data_3_12_to_3_13),
  .b_data_in(b_data_2_13_to_3_13),
  .c_data(c_data_3_13),
  .a_data_out(a_data_3_13_to_3_14),
  .b_data_out(b_data_3_13_to_4_13),
  .a_addr(a_addr_3_13_NC),
  .b_addr(b_addr_3_13_NC),
  .c_addr(c_addr_3_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 3_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_14_to_3_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_14_to_4_14;
  wire [`AWIDTH-1:0] a_addr_3_14_NC;
  wire [`AWIDTH-1:0] b_addr_3_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_14),
  .a_data(a_data_3_14_NC),
  .b_data(b_data_3_14_NC),
  .a_data_in(a_data_3_13_to_3_14),
  .b_data_in(b_data_2_14_to_3_14),
  .c_data(c_data_3_14),
  .a_data_out(a_data_3_14_to_3_15),
  .b_data_out(b_data_3_14_to_4_14),
  .a_addr(a_addr_3_14_NC),
  .b_addr(b_addr_3_14_NC),
  .c_addr(c_addr_3_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 3_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_15_to_3_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_15_to_4_15;
  wire [`AWIDTH-1:0] a_addr_3_15_NC;
  wire [`AWIDTH-1:0] b_addr_3_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_3_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_3_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_3_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_3_15),
  .a_data(a_data_3_15_NC),
  .b_data(b_data_3_15_NC),
  .a_data_in(a_data_3_14_to_3_15),
  .b_data_in(b_data_2_15_to_3_15),
  .c_data(c_data_3_15),
  .a_data_out(a_data_3_15_to_3_16),
  .b_data_out(b_data_3_15_to_4_15),
  .a_addr(a_addr_3_15_NC),
  .b_addr(b_addr_3_15_NC),
  .c_addr(c_addr_3_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd3),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 4_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_0_to_4_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_0_to_5_0;
  wire [`AWIDTH-1:0] b_addr_4_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_4_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_0),
  .a_data(a_data_4_0),
  .b_data(b_data_4_0_NC),
  .a_data_in(a_data_in_4_0_NC),
  .b_data_in(b_data_3_0_to_4_0),
  .c_data(c_data_4_0),
  .a_data_out(a_data_4_0_to_4_1),
  .b_data_out(b_data_4_0_to_5_0),
  .a_addr(a_addr_4_0),
  .b_addr(b_addr_4_0_NC),
  .c_addr(c_addr_4_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 4_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_1_to_4_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_1_to_5_1;
  wire [`AWIDTH-1:0] a_addr_4_1_NC;
  wire [`AWIDTH-1:0] b_addr_4_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_1),
  .a_data(a_data_4_1_NC),
  .b_data(b_data_4_1_NC),
  .a_data_in(a_data_4_0_to_4_1),
  .b_data_in(b_data_3_1_to_4_1),
  .c_data(c_data_4_1),
  .a_data_out(a_data_4_1_to_4_2),
  .b_data_out(b_data_4_1_to_5_1),
  .a_addr(a_addr_4_1_NC),
  .b_addr(b_addr_4_1_NC),
  .c_addr(c_addr_4_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 4_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_2_to_4_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_2_to_5_2;
  wire [`AWIDTH-1:0] a_addr_4_2_NC;
  wire [`AWIDTH-1:0] b_addr_4_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_2),
  .a_data(a_data_4_2_NC),
  .b_data(b_data_4_2_NC),
  .a_data_in(a_data_4_1_to_4_2),
  .b_data_in(b_data_3_2_to_4_2),
  .c_data(c_data_4_2),
  .a_data_out(a_data_4_2_to_4_3),
  .b_data_out(b_data_4_2_to_5_2),
  .a_addr(a_addr_4_2_NC),
  .b_addr(b_addr_4_2_NC),
  .c_addr(c_addr_4_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 4_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_3_to_4_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_3_to_5_3;
  wire [`AWIDTH-1:0] a_addr_4_3_NC;
  wire [`AWIDTH-1:0] b_addr_4_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_3),
  .a_data(a_data_4_3_NC),
  .b_data(b_data_4_3_NC),
  .a_data_in(a_data_4_2_to_4_3),
  .b_data_in(b_data_3_3_to_4_3),
  .c_data(c_data_4_3),
  .a_data_out(a_data_4_3_to_4_4),
  .b_data_out(b_data_4_3_to_5_3),
  .a_addr(a_addr_4_3_NC),
  .b_addr(b_addr_4_3_NC),
  .c_addr(c_addr_4_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 4_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_4_to_4_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_4_to_5_4;
  wire [`AWIDTH-1:0] a_addr_4_4_NC;
  wire [`AWIDTH-1:0] b_addr_4_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_4),
  .a_data(a_data_4_4_NC),
  .b_data(b_data_4_4_NC),
  .a_data_in(a_data_4_3_to_4_4),
  .b_data_in(b_data_3_4_to_4_4),
  .c_data(c_data_4_4),
  .a_data_out(a_data_4_4_to_4_5),
  .b_data_out(b_data_4_4_to_5_4),
  .a_addr(a_addr_4_4_NC),
  .b_addr(b_addr_4_4_NC),
  .c_addr(c_addr_4_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 4_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_5_to_4_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_5_to_5_5;
  wire [`AWIDTH-1:0] a_addr_4_5_NC;
  wire [`AWIDTH-1:0] b_addr_4_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_5),
  .a_data(a_data_4_5_NC),
  .b_data(b_data_4_5_NC),
  .a_data_in(a_data_4_4_to_4_5),
  .b_data_in(b_data_3_5_to_4_5),
  .c_data(c_data_4_5),
  .a_data_out(a_data_4_5_to_4_6),
  .b_data_out(b_data_4_5_to_5_5),
  .a_addr(a_addr_4_5_NC),
  .b_addr(b_addr_4_5_NC),
  .c_addr(c_addr_4_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 4_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_6_to_4_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_6_to_5_6;
  wire [`AWIDTH-1:0] a_addr_4_6_NC;
  wire [`AWIDTH-1:0] b_addr_4_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_6),
  .a_data(a_data_4_6_NC),
  .b_data(b_data_4_6_NC),
  .a_data_in(a_data_4_5_to_4_6),
  .b_data_in(b_data_3_6_to_4_6),
  .c_data(c_data_4_6),
  .a_data_out(a_data_4_6_to_4_7),
  .b_data_out(b_data_4_6_to_5_6),
  .a_addr(a_addr_4_6_NC),
  .b_addr(b_addr_4_6_NC),
  .c_addr(c_addr_4_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 4_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_7_to_4_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_7_to_5_7;
  wire [`AWIDTH-1:0] a_addr_4_7_NC;
  wire [`AWIDTH-1:0] b_addr_4_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_7),
  .a_data(a_data_4_7_NC),
  .b_data(b_data_4_7_NC),
  .a_data_in(a_data_4_6_to_4_7),
  .b_data_in(b_data_3_7_to_4_7),
  .c_data(c_data_4_7),
  .a_data_out(a_data_4_7_to_4_8),
  .b_data_out(b_data_4_7_to_5_7),
  .a_addr(a_addr_4_7_NC),
  .b_addr(b_addr_4_7_NC),
  .c_addr(c_addr_4_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 4_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_8_to_4_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_8_to_5_8;
  wire [`AWIDTH-1:0] a_addr_4_8_NC;
  wire [`AWIDTH-1:0] b_addr_4_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_8),
  .a_data(a_data_4_8_NC),
  .b_data(b_data_4_8_NC),
  .a_data_in(a_data_4_7_to_4_8),
  .b_data_in(b_data_3_8_to_4_8),
  .c_data(c_data_4_8),
  .a_data_out(a_data_4_8_to_4_9),
  .b_data_out(b_data_4_8_to_5_8),
  .a_addr(a_addr_4_8_NC),
  .b_addr(b_addr_4_8_NC),
  .c_addr(c_addr_4_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 4_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_9_to_4_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_9_to_5_9;
  wire [`AWIDTH-1:0] a_addr_4_9_NC;
  wire [`AWIDTH-1:0] b_addr_4_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_9),
  .a_data(a_data_4_9_NC),
  .b_data(b_data_4_9_NC),
  .a_data_in(a_data_4_8_to_4_9),
  .b_data_in(b_data_3_9_to_4_9),
  .c_data(c_data_4_9),
  .a_data_out(a_data_4_9_to_4_10),
  .b_data_out(b_data_4_9_to_5_9),
  .a_addr(a_addr_4_9_NC),
  .b_addr(b_addr_4_9_NC),
  .c_addr(c_addr_4_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 4_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_10_to_4_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_10_to_5_10;
  wire [`AWIDTH-1:0] a_addr_4_10_NC;
  wire [`AWIDTH-1:0] b_addr_4_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_10),
  .a_data(a_data_4_10_NC),
  .b_data(b_data_4_10_NC),
  .a_data_in(a_data_4_9_to_4_10),
  .b_data_in(b_data_3_10_to_4_10),
  .c_data(c_data_4_10),
  .a_data_out(a_data_4_10_to_4_11),
  .b_data_out(b_data_4_10_to_5_10),
  .a_addr(a_addr_4_10_NC),
  .b_addr(b_addr_4_10_NC),
  .c_addr(c_addr_4_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 4_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_11_to_4_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_11_to_5_11;
  wire [`AWIDTH-1:0] a_addr_4_11_NC;
  wire [`AWIDTH-1:0] b_addr_4_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_11),
  .a_data(a_data_4_11_NC),
  .b_data(b_data_4_11_NC),
  .a_data_in(a_data_4_10_to_4_11),
  .b_data_in(b_data_3_11_to_4_11),
  .c_data(c_data_4_11),
  .a_data_out(a_data_4_11_to_4_12),
  .b_data_out(b_data_4_11_to_5_11),
  .a_addr(a_addr_4_11_NC),
  .b_addr(b_addr_4_11_NC),
  .c_addr(c_addr_4_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 4_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_12_to_4_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_12_to_5_12;
  wire [`AWIDTH-1:0] a_addr_4_12_NC;
  wire [`AWIDTH-1:0] b_addr_4_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_12),
  .a_data(a_data_4_12_NC),
  .b_data(b_data_4_12_NC),
  .a_data_in(a_data_4_11_to_4_12),
  .b_data_in(b_data_3_12_to_4_12),
  .c_data(c_data_4_12),
  .a_data_out(a_data_4_12_to_4_13),
  .b_data_out(b_data_4_12_to_5_12),
  .a_addr(a_addr_4_12_NC),
  .b_addr(b_addr_4_12_NC),
  .c_addr(c_addr_4_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 4_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_13_to_4_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_13_to_5_13;
  wire [`AWIDTH-1:0] a_addr_4_13_NC;
  wire [`AWIDTH-1:0] b_addr_4_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_13),
  .a_data(a_data_4_13_NC),
  .b_data(b_data_4_13_NC),
  .a_data_in(a_data_4_12_to_4_13),
  .b_data_in(b_data_3_13_to_4_13),
  .c_data(c_data_4_13),
  .a_data_out(a_data_4_13_to_4_14),
  .b_data_out(b_data_4_13_to_5_13),
  .a_addr(a_addr_4_13_NC),
  .b_addr(b_addr_4_13_NC),
  .c_addr(c_addr_4_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 4_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_14_to_4_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_14_to_5_14;
  wire [`AWIDTH-1:0] a_addr_4_14_NC;
  wire [`AWIDTH-1:0] b_addr_4_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_14),
  .a_data(a_data_4_14_NC),
  .b_data(b_data_4_14_NC),
  .a_data_in(a_data_4_13_to_4_14),
  .b_data_in(b_data_3_14_to_4_14),
  .c_data(c_data_4_14),
  .a_data_out(a_data_4_14_to_4_15),
  .b_data_out(b_data_4_14_to_5_14),
  .a_addr(a_addr_4_14_NC),
  .b_addr(b_addr_4_14_NC),
  .c_addr(c_addr_4_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 4_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_15_to_4_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_15_to_5_15;
  wire [`AWIDTH-1:0] a_addr_4_15_NC;
  wire [`AWIDTH-1:0] b_addr_4_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_4_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_4_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_4_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_4_15),
  .a_data(a_data_4_15_NC),
  .b_data(b_data_4_15_NC),
  .a_data_in(a_data_4_14_to_4_15),
  .b_data_in(b_data_3_15_to_4_15),
  .c_data(c_data_4_15),
  .a_data_out(a_data_4_15_to_4_16),
  .b_data_out(b_data_4_15_to_5_15),
  .a_addr(a_addr_4_15_NC),
  .b_addr(b_addr_4_15_NC),
  .c_addr(c_addr_4_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd4),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 5_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_0_to_5_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_0_to_6_0;
  wire [`AWIDTH-1:0] b_addr_5_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_5_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_0),
  .a_data(a_data_5_0),
  .b_data(b_data_5_0_NC),
  .a_data_in(a_data_in_5_0_NC),
  .b_data_in(b_data_4_0_to_5_0),
  .c_data(c_data_5_0),
  .a_data_out(a_data_5_0_to_5_1),
  .b_data_out(b_data_5_0_to_6_0),
  .a_addr(a_addr_5_0),
  .b_addr(b_addr_5_0_NC),
  .c_addr(c_addr_5_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 5_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_1_to_5_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_1_to_6_1;
  wire [`AWIDTH-1:0] a_addr_5_1_NC;
  wire [`AWIDTH-1:0] b_addr_5_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_1),
  .a_data(a_data_5_1_NC),
  .b_data(b_data_5_1_NC),
  .a_data_in(a_data_5_0_to_5_1),
  .b_data_in(b_data_4_1_to_5_1),
  .c_data(c_data_5_1),
  .a_data_out(a_data_5_1_to_5_2),
  .b_data_out(b_data_5_1_to_6_1),
  .a_addr(a_addr_5_1_NC),
  .b_addr(b_addr_5_1_NC),
  .c_addr(c_addr_5_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 5_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_2_to_5_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_2_to_6_2;
  wire [`AWIDTH-1:0] a_addr_5_2_NC;
  wire [`AWIDTH-1:0] b_addr_5_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_2),
  .a_data(a_data_5_2_NC),
  .b_data(b_data_5_2_NC),
  .a_data_in(a_data_5_1_to_5_2),
  .b_data_in(b_data_4_2_to_5_2),
  .c_data(c_data_5_2),
  .a_data_out(a_data_5_2_to_5_3),
  .b_data_out(b_data_5_2_to_6_2),
  .a_addr(a_addr_5_2_NC),
  .b_addr(b_addr_5_2_NC),
  .c_addr(c_addr_5_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 5_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_3_to_5_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_3_to_6_3;
  wire [`AWIDTH-1:0] a_addr_5_3_NC;
  wire [`AWIDTH-1:0] b_addr_5_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_3),
  .a_data(a_data_5_3_NC),
  .b_data(b_data_5_3_NC),
  .a_data_in(a_data_5_2_to_5_3),
  .b_data_in(b_data_4_3_to_5_3),
  .c_data(c_data_5_3),
  .a_data_out(a_data_5_3_to_5_4),
  .b_data_out(b_data_5_3_to_6_3),
  .a_addr(a_addr_5_3_NC),
  .b_addr(b_addr_5_3_NC),
  .c_addr(c_addr_5_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 5_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_4_to_5_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_4_to_6_4;
  wire [`AWIDTH-1:0] a_addr_5_4_NC;
  wire [`AWIDTH-1:0] b_addr_5_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_4),
  .a_data(a_data_5_4_NC),
  .b_data(b_data_5_4_NC),
  .a_data_in(a_data_5_3_to_5_4),
  .b_data_in(b_data_4_4_to_5_4),
  .c_data(c_data_5_4),
  .a_data_out(a_data_5_4_to_5_5),
  .b_data_out(b_data_5_4_to_6_4),
  .a_addr(a_addr_5_4_NC),
  .b_addr(b_addr_5_4_NC),
  .c_addr(c_addr_5_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 5_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_5_to_5_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_5_to_6_5;
  wire [`AWIDTH-1:0] a_addr_5_5_NC;
  wire [`AWIDTH-1:0] b_addr_5_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_5),
  .a_data(a_data_5_5_NC),
  .b_data(b_data_5_5_NC),
  .a_data_in(a_data_5_4_to_5_5),
  .b_data_in(b_data_4_5_to_5_5),
  .c_data(c_data_5_5),
  .a_data_out(a_data_5_5_to_5_6),
  .b_data_out(b_data_5_5_to_6_5),
  .a_addr(a_addr_5_5_NC),
  .b_addr(b_addr_5_5_NC),
  .c_addr(c_addr_5_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 5_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_6_to_5_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_6_to_6_6;
  wire [`AWIDTH-1:0] a_addr_5_6_NC;
  wire [`AWIDTH-1:0] b_addr_5_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_6),
  .a_data(a_data_5_6_NC),
  .b_data(b_data_5_6_NC),
  .a_data_in(a_data_5_5_to_5_6),
  .b_data_in(b_data_4_6_to_5_6),
  .c_data(c_data_5_6),
  .a_data_out(a_data_5_6_to_5_7),
  .b_data_out(b_data_5_6_to_6_6),
  .a_addr(a_addr_5_6_NC),
  .b_addr(b_addr_5_6_NC),
  .c_addr(c_addr_5_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 5_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_7_to_5_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_7_to_6_7;
  wire [`AWIDTH-1:0] a_addr_5_7_NC;
  wire [`AWIDTH-1:0] b_addr_5_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_7),
  .a_data(a_data_5_7_NC),
  .b_data(b_data_5_7_NC),
  .a_data_in(a_data_5_6_to_5_7),
  .b_data_in(b_data_4_7_to_5_7),
  .c_data(c_data_5_7),
  .a_data_out(a_data_5_7_to_5_8),
  .b_data_out(b_data_5_7_to_6_7),
  .a_addr(a_addr_5_7_NC),
  .b_addr(b_addr_5_7_NC),
  .c_addr(c_addr_5_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 5_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_8_to_5_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_8_to_6_8;
  wire [`AWIDTH-1:0] a_addr_5_8_NC;
  wire [`AWIDTH-1:0] b_addr_5_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_8),
  .a_data(a_data_5_8_NC),
  .b_data(b_data_5_8_NC),
  .a_data_in(a_data_5_7_to_5_8),
  .b_data_in(b_data_4_8_to_5_8),
  .c_data(c_data_5_8),
  .a_data_out(a_data_5_8_to_5_9),
  .b_data_out(b_data_5_8_to_6_8),
  .a_addr(a_addr_5_8_NC),
  .b_addr(b_addr_5_8_NC),
  .c_addr(c_addr_5_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 5_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_9_to_5_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_9_to_6_9;
  wire [`AWIDTH-1:0] a_addr_5_9_NC;
  wire [`AWIDTH-1:0] b_addr_5_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_9),
  .a_data(a_data_5_9_NC),
  .b_data(b_data_5_9_NC),
  .a_data_in(a_data_5_8_to_5_9),
  .b_data_in(b_data_4_9_to_5_9),
  .c_data(c_data_5_9),
  .a_data_out(a_data_5_9_to_5_10),
  .b_data_out(b_data_5_9_to_6_9),
  .a_addr(a_addr_5_9_NC),
  .b_addr(b_addr_5_9_NC),
  .c_addr(c_addr_5_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 5_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_10_to_5_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_10_to_6_10;
  wire [`AWIDTH-1:0] a_addr_5_10_NC;
  wire [`AWIDTH-1:0] b_addr_5_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_10),
  .a_data(a_data_5_10_NC),
  .b_data(b_data_5_10_NC),
  .a_data_in(a_data_5_9_to_5_10),
  .b_data_in(b_data_4_10_to_5_10),
  .c_data(c_data_5_10),
  .a_data_out(a_data_5_10_to_5_11),
  .b_data_out(b_data_5_10_to_6_10),
  .a_addr(a_addr_5_10_NC),
  .b_addr(b_addr_5_10_NC),
  .c_addr(c_addr_5_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 5_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_11_to_5_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_11_to_6_11;
  wire [`AWIDTH-1:0] a_addr_5_11_NC;
  wire [`AWIDTH-1:0] b_addr_5_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_11),
  .a_data(a_data_5_11_NC),
  .b_data(b_data_5_11_NC),
  .a_data_in(a_data_5_10_to_5_11),
  .b_data_in(b_data_4_11_to_5_11),
  .c_data(c_data_5_11),
  .a_data_out(a_data_5_11_to_5_12),
  .b_data_out(b_data_5_11_to_6_11),
  .a_addr(a_addr_5_11_NC),
  .b_addr(b_addr_5_11_NC),
  .c_addr(c_addr_5_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 5_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_12_to_5_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_12_to_6_12;
  wire [`AWIDTH-1:0] a_addr_5_12_NC;
  wire [`AWIDTH-1:0] b_addr_5_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_12),
  .a_data(a_data_5_12_NC),
  .b_data(b_data_5_12_NC),
  .a_data_in(a_data_5_11_to_5_12),
  .b_data_in(b_data_4_12_to_5_12),
  .c_data(c_data_5_12),
  .a_data_out(a_data_5_12_to_5_13),
  .b_data_out(b_data_5_12_to_6_12),
  .a_addr(a_addr_5_12_NC),
  .b_addr(b_addr_5_12_NC),
  .c_addr(c_addr_5_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 5_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_13_to_5_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_13_to_6_13;
  wire [`AWIDTH-1:0] a_addr_5_13_NC;
  wire [`AWIDTH-1:0] b_addr_5_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_13),
  .a_data(a_data_5_13_NC),
  .b_data(b_data_5_13_NC),
  .a_data_in(a_data_5_12_to_5_13),
  .b_data_in(b_data_4_13_to_5_13),
  .c_data(c_data_5_13),
  .a_data_out(a_data_5_13_to_5_14),
  .b_data_out(b_data_5_13_to_6_13),
  .a_addr(a_addr_5_13_NC),
  .b_addr(b_addr_5_13_NC),
  .c_addr(c_addr_5_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 5_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_14_to_5_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_14_to_6_14;
  wire [`AWIDTH-1:0] a_addr_5_14_NC;
  wire [`AWIDTH-1:0] b_addr_5_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_14),
  .a_data(a_data_5_14_NC),
  .b_data(b_data_5_14_NC),
  .a_data_in(a_data_5_13_to_5_14),
  .b_data_in(b_data_4_14_to_5_14),
  .c_data(c_data_5_14),
  .a_data_out(a_data_5_14_to_5_15),
  .b_data_out(b_data_5_14_to_6_14),
  .a_addr(a_addr_5_14_NC),
  .b_addr(b_addr_5_14_NC),
  .c_addr(c_addr_5_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 5_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_15_to_5_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_15_to_6_15;
  wire [`AWIDTH-1:0] a_addr_5_15_NC;
  wire [`AWIDTH-1:0] b_addr_5_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_5_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_5_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_5_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_5_15),
  .a_data(a_data_5_15_NC),
  .b_data(b_data_5_15_NC),
  .a_data_in(a_data_5_14_to_5_15),
  .b_data_in(b_data_4_15_to_5_15),
  .c_data(c_data_5_15),
  .a_data_out(a_data_5_15_to_5_16),
  .b_data_out(b_data_5_15_to_6_15),
  .a_addr(a_addr_5_15_NC),
  .b_addr(b_addr_5_15_NC),
  .c_addr(c_addr_5_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd5),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 6_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_0_to_6_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_0_to_7_0;
  wire [`AWIDTH-1:0] b_addr_6_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_6_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_0),
  .a_data(a_data_6_0),
  .b_data(b_data_6_0_NC),
  .a_data_in(a_data_in_6_0_NC),
  .b_data_in(b_data_5_0_to_6_0),
  .c_data(c_data_6_0),
  .a_data_out(a_data_6_0_to_6_1),
  .b_data_out(b_data_6_0_to_7_0),
  .a_addr(a_addr_6_0),
  .b_addr(b_addr_6_0_NC),
  .c_addr(c_addr_6_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 6_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_1_to_6_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_1_to_7_1;
  wire [`AWIDTH-1:0] a_addr_6_1_NC;
  wire [`AWIDTH-1:0] b_addr_6_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_1),
  .a_data(a_data_6_1_NC),
  .b_data(b_data_6_1_NC),
  .a_data_in(a_data_6_0_to_6_1),
  .b_data_in(b_data_5_1_to_6_1),
  .c_data(c_data_6_1),
  .a_data_out(a_data_6_1_to_6_2),
  .b_data_out(b_data_6_1_to_7_1),
  .a_addr(a_addr_6_1_NC),
  .b_addr(b_addr_6_1_NC),
  .c_addr(c_addr_6_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 6_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_2_to_6_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_2_to_7_2;
  wire [`AWIDTH-1:0] a_addr_6_2_NC;
  wire [`AWIDTH-1:0] b_addr_6_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_2),
  .a_data(a_data_6_2_NC),
  .b_data(b_data_6_2_NC),
  .a_data_in(a_data_6_1_to_6_2),
  .b_data_in(b_data_5_2_to_6_2),
  .c_data(c_data_6_2),
  .a_data_out(a_data_6_2_to_6_3),
  .b_data_out(b_data_6_2_to_7_2),
  .a_addr(a_addr_6_2_NC),
  .b_addr(b_addr_6_2_NC),
  .c_addr(c_addr_6_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 6_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_3_to_6_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_3_to_7_3;
  wire [`AWIDTH-1:0] a_addr_6_3_NC;
  wire [`AWIDTH-1:0] b_addr_6_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_3),
  .a_data(a_data_6_3_NC),
  .b_data(b_data_6_3_NC),
  .a_data_in(a_data_6_2_to_6_3),
  .b_data_in(b_data_5_3_to_6_3),
  .c_data(c_data_6_3),
  .a_data_out(a_data_6_3_to_6_4),
  .b_data_out(b_data_6_3_to_7_3),
  .a_addr(a_addr_6_3_NC),
  .b_addr(b_addr_6_3_NC),
  .c_addr(c_addr_6_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 6_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_4_to_6_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_4_to_7_4;
  wire [`AWIDTH-1:0] a_addr_6_4_NC;
  wire [`AWIDTH-1:0] b_addr_6_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_4),
  .a_data(a_data_6_4_NC),
  .b_data(b_data_6_4_NC),
  .a_data_in(a_data_6_3_to_6_4),
  .b_data_in(b_data_5_4_to_6_4),
  .c_data(c_data_6_4),
  .a_data_out(a_data_6_4_to_6_5),
  .b_data_out(b_data_6_4_to_7_4),
  .a_addr(a_addr_6_4_NC),
  .b_addr(b_addr_6_4_NC),
  .c_addr(c_addr_6_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 6_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_5_to_6_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_5_to_7_5;
  wire [`AWIDTH-1:0] a_addr_6_5_NC;
  wire [`AWIDTH-1:0] b_addr_6_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_5),
  .a_data(a_data_6_5_NC),
  .b_data(b_data_6_5_NC),
  .a_data_in(a_data_6_4_to_6_5),
  .b_data_in(b_data_5_5_to_6_5),
  .c_data(c_data_6_5),
  .a_data_out(a_data_6_5_to_6_6),
  .b_data_out(b_data_6_5_to_7_5),
  .a_addr(a_addr_6_5_NC),
  .b_addr(b_addr_6_5_NC),
  .c_addr(c_addr_6_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 6_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_6_to_6_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_6_to_7_6;
  wire [`AWIDTH-1:0] a_addr_6_6_NC;
  wire [`AWIDTH-1:0] b_addr_6_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_6),
  .a_data(a_data_6_6_NC),
  .b_data(b_data_6_6_NC),
  .a_data_in(a_data_6_5_to_6_6),
  .b_data_in(b_data_5_6_to_6_6),
  .c_data(c_data_6_6),
  .a_data_out(a_data_6_6_to_6_7),
  .b_data_out(b_data_6_6_to_7_6),
  .a_addr(a_addr_6_6_NC),
  .b_addr(b_addr_6_6_NC),
  .c_addr(c_addr_6_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 6_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_7_to_6_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_7_to_7_7;
  wire [`AWIDTH-1:0] a_addr_6_7_NC;
  wire [`AWIDTH-1:0] b_addr_6_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_7),
  .a_data(a_data_6_7_NC),
  .b_data(b_data_6_7_NC),
  .a_data_in(a_data_6_6_to_6_7),
  .b_data_in(b_data_5_7_to_6_7),
  .c_data(c_data_6_7),
  .a_data_out(a_data_6_7_to_6_8),
  .b_data_out(b_data_6_7_to_7_7),
  .a_addr(a_addr_6_7_NC),
  .b_addr(b_addr_6_7_NC),
  .c_addr(c_addr_6_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 6_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_8_to_6_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_8_to_7_8;
  wire [`AWIDTH-1:0] a_addr_6_8_NC;
  wire [`AWIDTH-1:0] b_addr_6_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_8),
  .a_data(a_data_6_8_NC),
  .b_data(b_data_6_8_NC),
  .a_data_in(a_data_6_7_to_6_8),
  .b_data_in(b_data_5_8_to_6_8),
  .c_data(c_data_6_8),
  .a_data_out(a_data_6_8_to_6_9),
  .b_data_out(b_data_6_8_to_7_8),
  .a_addr(a_addr_6_8_NC),
  .b_addr(b_addr_6_8_NC),
  .c_addr(c_addr_6_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 6_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_9_to_6_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_9_to_7_9;
  wire [`AWIDTH-1:0] a_addr_6_9_NC;
  wire [`AWIDTH-1:0] b_addr_6_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_9),
  .a_data(a_data_6_9_NC),
  .b_data(b_data_6_9_NC),
  .a_data_in(a_data_6_8_to_6_9),
  .b_data_in(b_data_5_9_to_6_9),
  .c_data(c_data_6_9),
  .a_data_out(a_data_6_9_to_6_10),
  .b_data_out(b_data_6_9_to_7_9),
  .a_addr(a_addr_6_9_NC),
  .b_addr(b_addr_6_9_NC),
  .c_addr(c_addr_6_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 6_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_10_to_6_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_10_to_7_10;
  wire [`AWIDTH-1:0] a_addr_6_10_NC;
  wire [`AWIDTH-1:0] b_addr_6_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_10),
  .a_data(a_data_6_10_NC),
  .b_data(b_data_6_10_NC),
  .a_data_in(a_data_6_9_to_6_10),
  .b_data_in(b_data_5_10_to_6_10),
  .c_data(c_data_6_10),
  .a_data_out(a_data_6_10_to_6_11),
  .b_data_out(b_data_6_10_to_7_10),
  .a_addr(a_addr_6_10_NC),
  .b_addr(b_addr_6_10_NC),
  .c_addr(c_addr_6_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 6_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_11_to_6_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_11_to_7_11;
  wire [`AWIDTH-1:0] a_addr_6_11_NC;
  wire [`AWIDTH-1:0] b_addr_6_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_11),
  .a_data(a_data_6_11_NC),
  .b_data(b_data_6_11_NC),
  .a_data_in(a_data_6_10_to_6_11),
  .b_data_in(b_data_5_11_to_6_11),
  .c_data(c_data_6_11),
  .a_data_out(a_data_6_11_to_6_12),
  .b_data_out(b_data_6_11_to_7_11),
  .a_addr(a_addr_6_11_NC),
  .b_addr(b_addr_6_11_NC),
  .c_addr(c_addr_6_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 6_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_12_to_6_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_12_to_7_12;
  wire [`AWIDTH-1:0] a_addr_6_12_NC;
  wire [`AWIDTH-1:0] b_addr_6_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_12),
  .a_data(a_data_6_12_NC),
  .b_data(b_data_6_12_NC),
  .a_data_in(a_data_6_11_to_6_12),
  .b_data_in(b_data_5_12_to_6_12),
  .c_data(c_data_6_12),
  .a_data_out(a_data_6_12_to_6_13),
  .b_data_out(b_data_6_12_to_7_12),
  .a_addr(a_addr_6_12_NC),
  .b_addr(b_addr_6_12_NC),
  .c_addr(c_addr_6_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 6_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_13_to_6_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_13_to_7_13;
  wire [`AWIDTH-1:0] a_addr_6_13_NC;
  wire [`AWIDTH-1:0] b_addr_6_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_13),
  .a_data(a_data_6_13_NC),
  .b_data(b_data_6_13_NC),
  .a_data_in(a_data_6_12_to_6_13),
  .b_data_in(b_data_5_13_to_6_13),
  .c_data(c_data_6_13),
  .a_data_out(a_data_6_13_to_6_14),
  .b_data_out(b_data_6_13_to_7_13),
  .a_addr(a_addr_6_13_NC),
  .b_addr(b_addr_6_13_NC),
  .c_addr(c_addr_6_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 6_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_14_to_6_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_14_to_7_14;
  wire [`AWIDTH-1:0] a_addr_6_14_NC;
  wire [`AWIDTH-1:0] b_addr_6_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_14),
  .a_data(a_data_6_14_NC),
  .b_data(b_data_6_14_NC),
  .a_data_in(a_data_6_13_to_6_14),
  .b_data_in(b_data_5_14_to_6_14),
  .c_data(c_data_6_14),
  .a_data_out(a_data_6_14_to_6_15),
  .b_data_out(b_data_6_14_to_7_14),
  .a_addr(a_addr_6_14_NC),
  .b_addr(b_addr_6_14_NC),
  .c_addr(c_addr_6_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 6_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_15_to_6_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_15_to_7_15;
  wire [`AWIDTH-1:0] a_addr_6_15_NC;
  wire [`AWIDTH-1:0] b_addr_6_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_6_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_6_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_6_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_6_15),
  .a_data(a_data_6_15_NC),
  .b_data(b_data_6_15_NC),
  .a_data_in(a_data_6_14_to_6_15),
  .b_data_in(b_data_5_15_to_6_15),
  .c_data(c_data_6_15),
  .a_data_out(a_data_6_15_to_6_16),
  .b_data_out(b_data_6_15_to_7_15),
  .a_addr(a_addr_6_15_NC),
  .b_addr(b_addr_6_15_NC),
  .c_addr(c_addr_6_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd6),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 7_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_0_to_7_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_0_to_8_0;
  wire [`AWIDTH-1:0] b_addr_7_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_7_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_0),
  .a_data(a_data_7_0),
  .b_data(b_data_7_0_NC),
  .a_data_in(a_data_in_7_0_NC),
  .b_data_in(b_data_6_0_to_7_0),
  .c_data(c_data_7_0),
  .a_data_out(a_data_7_0_to_7_1),
  .b_data_out(b_data_7_0_to_8_0),
  .a_addr(a_addr_7_0),
  .b_addr(b_addr_7_0_NC),
  .c_addr(c_addr_7_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 7_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_1_to_7_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_1_to_8_1;
  wire [`AWIDTH-1:0] a_addr_7_1_NC;
  wire [`AWIDTH-1:0] b_addr_7_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_1),
  .a_data(a_data_7_1_NC),
  .b_data(b_data_7_1_NC),
  .a_data_in(a_data_7_0_to_7_1),
  .b_data_in(b_data_6_1_to_7_1),
  .c_data(c_data_7_1),
  .a_data_out(a_data_7_1_to_7_2),
  .b_data_out(b_data_7_1_to_8_1),
  .a_addr(a_addr_7_1_NC),
  .b_addr(b_addr_7_1_NC),
  .c_addr(c_addr_7_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 7_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_2_to_7_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_2_to_8_2;
  wire [`AWIDTH-1:0] a_addr_7_2_NC;
  wire [`AWIDTH-1:0] b_addr_7_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_2),
  .a_data(a_data_7_2_NC),
  .b_data(b_data_7_2_NC),
  .a_data_in(a_data_7_1_to_7_2),
  .b_data_in(b_data_6_2_to_7_2),
  .c_data(c_data_7_2),
  .a_data_out(a_data_7_2_to_7_3),
  .b_data_out(b_data_7_2_to_8_2),
  .a_addr(a_addr_7_2_NC),
  .b_addr(b_addr_7_2_NC),
  .c_addr(c_addr_7_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 7_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_3_to_7_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_3_to_8_3;
  wire [`AWIDTH-1:0] a_addr_7_3_NC;
  wire [`AWIDTH-1:0] b_addr_7_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_3),
  .a_data(a_data_7_3_NC),
  .b_data(b_data_7_3_NC),
  .a_data_in(a_data_7_2_to_7_3),
  .b_data_in(b_data_6_3_to_7_3),
  .c_data(c_data_7_3),
  .a_data_out(a_data_7_3_to_7_4),
  .b_data_out(b_data_7_3_to_8_3),
  .a_addr(a_addr_7_3_NC),
  .b_addr(b_addr_7_3_NC),
  .c_addr(c_addr_7_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 7_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_4_to_7_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_4_to_8_4;
  wire [`AWIDTH-1:0] a_addr_7_4_NC;
  wire [`AWIDTH-1:0] b_addr_7_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_4),
  .a_data(a_data_7_4_NC),
  .b_data(b_data_7_4_NC),
  .a_data_in(a_data_7_3_to_7_4),
  .b_data_in(b_data_6_4_to_7_4),
  .c_data(c_data_7_4),
  .a_data_out(a_data_7_4_to_7_5),
  .b_data_out(b_data_7_4_to_8_4),
  .a_addr(a_addr_7_4_NC),
  .b_addr(b_addr_7_4_NC),
  .c_addr(c_addr_7_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 7_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_5_to_7_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_5_to_8_5;
  wire [`AWIDTH-1:0] a_addr_7_5_NC;
  wire [`AWIDTH-1:0] b_addr_7_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_5),
  .a_data(a_data_7_5_NC),
  .b_data(b_data_7_5_NC),
  .a_data_in(a_data_7_4_to_7_5),
  .b_data_in(b_data_6_5_to_7_5),
  .c_data(c_data_7_5),
  .a_data_out(a_data_7_5_to_7_6),
  .b_data_out(b_data_7_5_to_8_5),
  .a_addr(a_addr_7_5_NC),
  .b_addr(b_addr_7_5_NC),
  .c_addr(c_addr_7_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 7_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_6_to_7_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_6_to_8_6;
  wire [`AWIDTH-1:0] a_addr_7_6_NC;
  wire [`AWIDTH-1:0] b_addr_7_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_6),
  .a_data(a_data_7_6_NC),
  .b_data(b_data_7_6_NC),
  .a_data_in(a_data_7_5_to_7_6),
  .b_data_in(b_data_6_6_to_7_6),
  .c_data(c_data_7_6),
  .a_data_out(a_data_7_6_to_7_7),
  .b_data_out(b_data_7_6_to_8_6),
  .a_addr(a_addr_7_6_NC),
  .b_addr(b_addr_7_6_NC),
  .c_addr(c_addr_7_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 7_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_7_to_7_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_7_to_8_7;
  wire [`AWIDTH-1:0] a_addr_7_7_NC;
  wire [`AWIDTH-1:0] b_addr_7_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_7),
  .a_data(a_data_7_7_NC),
  .b_data(b_data_7_7_NC),
  .a_data_in(a_data_7_6_to_7_7),
  .b_data_in(b_data_6_7_to_7_7),
  .c_data(c_data_7_7),
  .a_data_out(a_data_7_7_to_7_8),
  .b_data_out(b_data_7_7_to_8_7),
  .a_addr(a_addr_7_7_NC),
  .b_addr(b_addr_7_7_NC),
  .c_addr(c_addr_7_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 7_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_8_to_7_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_8_to_8_8;
  wire [`AWIDTH-1:0] a_addr_7_8_NC;
  wire [`AWIDTH-1:0] b_addr_7_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_8),
  .a_data(a_data_7_8_NC),
  .b_data(b_data_7_8_NC),
  .a_data_in(a_data_7_7_to_7_8),
  .b_data_in(b_data_6_8_to_7_8),
  .c_data(c_data_7_8),
  .a_data_out(a_data_7_8_to_7_9),
  .b_data_out(b_data_7_8_to_8_8),
  .a_addr(a_addr_7_8_NC),
  .b_addr(b_addr_7_8_NC),
  .c_addr(c_addr_7_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 7_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_9_to_7_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_9_to_8_9;
  wire [`AWIDTH-1:0] a_addr_7_9_NC;
  wire [`AWIDTH-1:0] b_addr_7_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_9),
  .a_data(a_data_7_9_NC),
  .b_data(b_data_7_9_NC),
  .a_data_in(a_data_7_8_to_7_9),
  .b_data_in(b_data_6_9_to_7_9),
  .c_data(c_data_7_9),
  .a_data_out(a_data_7_9_to_7_10),
  .b_data_out(b_data_7_9_to_8_9),
  .a_addr(a_addr_7_9_NC),
  .b_addr(b_addr_7_9_NC),
  .c_addr(c_addr_7_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 7_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_10_to_7_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_10_to_8_10;
  wire [`AWIDTH-1:0] a_addr_7_10_NC;
  wire [`AWIDTH-1:0] b_addr_7_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_10),
  .a_data(a_data_7_10_NC),
  .b_data(b_data_7_10_NC),
  .a_data_in(a_data_7_9_to_7_10),
  .b_data_in(b_data_6_10_to_7_10),
  .c_data(c_data_7_10),
  .a_data_out(a_data_7_10_to_7_11),
  .b_data_out(b_data_7_10_to_8_10),
  .a_addr(a_addr_7_10_NC),
  .b_addr(b_addr_7_10_NC),
  .c_addr(c_addr_7_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 7_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_11_to_7_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_11_to_8_11;
  wire [`AWIDTH-1:0] a_addr_7_11_NC;
  wire [`AWIDTH-1:0] b_addr_7_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_11),
  .a_data(a_data_7_11_NC),
  .b_data(b_data_7_11_NC),
  .a_data_in(a_data_7_10_to_7_11),
  .b_data_in(b_data_6_11_to_7_11),
  .c_data(c_data_7_11),
  .a_data_out(a_data_7_11_to_7_12),
  .b_data_out(b_data_7_11_to_8_11),
  .a_addr(a_addr_7_11_NC),
  .b_addr(b_addr_7_11_NC),
  .c_addr(c_addr_7_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 7_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_12_to_7_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_12_to_8_12;
  wire [`AWIDTH-1:0] a_addr_7_12_NC;
  wire [`AWIDTH-1:0] b_addr_7_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_12),
  .a_data(a_data_7_12_NC),
  .b_data(b_data_7_12_NC),
  .a_data_in(a_data_7_11_to_7_12),
  .b_data_in(b_data_6_12_to_7_12),
  .c_data(c_data_7_12),
  .a_data_out(a_data_7_12_to_7_13),
  .b_data_out(b_data_7_12_to_8_12),
  .a_addr(a_addr_7_12_NC),
  .b_addr(b_addr_7_12_NC),
  .c_addr(c_addr_7_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 7_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_13_to_7_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_13_to_8_13;
  wire [`AWIDTH-1:0] a_addr_7_13_NC;
  wire [`AWIDTH-1:0] b_addr_7_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_13),
  .a_data(a_data_7_13_NC),
  .b_data(b_data_7_13_NC),
  .a_data_in(a_data_7_12_to_7_13),
  .b_data_in(b_data_6_13_to_7_13),
  .c_data(c_data_7_13),
  .a_data_out(a_data_7_13_to_7_14),
  .b_data_out(b_data_7_13_to_8_13),
  .a_addr(a_addr_7_13_NC),
  .b_addr(b_addr_7_13_NC),
  .c_addr(c_addr_7_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 7_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_14_to_7_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_14_to_8_14;
  wire [`AWIDTH-1:0] a_addr_7_14_NC;
  wire [`AWIDTH-1:0] b_addr_7_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_14),
  .a_data(a_data_7_14_NC),
  .b_data(b_data_7_14_NC),
  .a_data_in(a_data_7_13_to_7_14),
  .b_data_in(b_data_6_14_to_7_14),
  .c_data(c_data_7_14),
  .a_data_out(a_data_7_14_to_7_15),
  .b_data_out(b_data_7_14_to_8_14),
  .a_addr(a_addr_7_14_NC),
  .b_addr(b_addr_7_14_NC),
  .c_addr(c_addr_7_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 7_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_15_to_7_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_15_to_8_15;
  wire [`AWIDTH-1:0] a_addr_7_15_NC;
  wire [`AWIDTH-1:0] b_addr_7_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_7_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_7_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_7_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_7_15),
  .a_data(a_data_7_15_NC),
  .b_data(b_data_7_15_NC),
  .a_data_in(a_data_7_14_to_7_15),
  .b_data_in(b_data_6_15_to_7_15),
  .c_data(c_data_7_15),
  .a_data_out(a_data_7_15_to_7_16),
  .b_data_out(b_data_7_15_to_8_15),
  .a_addr(a_addr_7_15_NC),
  .b_addr(b_addr_7_15_NC),
  .c_addr(c_addr_7_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd7),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 8_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_0_to_8_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_0_to_9_0;
  wire [`AWIDTH-1:0] b_addr_8_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_8_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_0),
  .a_data(a_data_8_0),
  .b_data(b_data_8_0_NC),
  .a_data_in(a_data_in_8_0_NC),
  .b_data_in(b_data_7_0_to_8_0),
  .c_data(c_data_8_0),
  .a_data_out(a_data_8_0_to_8_1),
  .b_data_out(b_data_8_0_to_9_0),
  .a_addr(a_addr_8_0),
  .b_addr(b_addr_8_0_NC),
  .c_addr(c_addr_8_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 8_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_1_to_8_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_1_to_9_1;
  wire [`AWIDTH-1:0] a_addr_8_1_NC;
  wire [`AWIDTH-1:0] b_addr_8_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_1),
  .a_data(a_data_8_1_NC),
  .b_data(b_data_8_1_NC),
  .a_data_in(a_data_8_0_to_8_1),
  .b_data_in(b_data_7_1_to_8_1),
  .c_data(c_data_8_1),
  .a_data_out(a_data_8_1_to_8_2),
  .b_data_out(b_data_8_1_to_9_1),
  .a_addr(a_addr_8_1_NC),
  .b_addr(b_addr_8_1_NC),
  .c_addr(c_addr_8_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 8_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_2_to_8_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_2_to_9_2;
  wire [`AWIDTH-1:0] a_addr_8_2_NC;
  wire [`AWIDTH-1:0] b_addr_8_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_2),
  .a_data(a_data_8_2_NC),
  .b_data(b_data_8_2_NC),
  .a_data_in(a_data_8_1_to_8_2),
  .b_data_in(b_data_7_2_to_8_2),
  .c_data(c_data_8_2),
  .a_data_out(a_data_8_2_to_8_3),
  .b_data_out(b_data_8_2_to_9_2),
  .a_addr(a_addr_8_2_NC),
  .b_addr(b_addr_8_2_NC),
  .c_addr(c_addr_8_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 8_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_3_to_8_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_3_to_9_3;
  wire [`AWIDTH-1:0] a_addr_8_3_NC;
  wire [`AWIDTH-1:0] b_addr_8_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_3),
  .a_data(a_data_8_3_NC),
  .b_data(b_data_8_3_NC),
  .a_data_in(a_data_8_2_to_8_3),
  .b_data_in(b_data_7_3_to_8_3),
  .c_data(c_data_8_3),
  .a_data_out(a_data_8_3_to_8_4),
  .b_data_out(b_data_8_3_to_9_3),
  .a_addr(a_addr_8_3_NC),
  .b_addr(b_addr_8_3_NC),
  .c_addr(c_addr_8_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 8_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_4_to_8_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_4_to_9_4;
  wire [`AWIDTH-1:0] a_addr_8_4_NC;
  wire [`AWIDTH-1:0] b_addr_8_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_4),
  .a_data(a_data_8_4_NC),
  .b_data(b_data_8_4_NC),
  .a_data_in(a_data_8_3_to_8_4),
  .b_data_in(b_data_7_4_to_8_4),
  .c_data(c_data_8_4),
  .a_data_out(a_data_8_4_to_8_5),
  .b_data_out(b_data_8_4_to_9_4),
  .a_addr(a_addr_8_4_NC),
  .b_addr(b_addr_8_4_NC),
  .c_addr(c_addr_8_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 8_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_5_to_8_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_5_to_9_5;
  wire [`AWIDTH-1:0] a_addr_8_5_NC;
  wire [`AWIDTH-1:0] b_addr_8_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_5),
  .a_data(a_data_8_5_NC),
  .b_data(b_data_8_5_NC),
  .a_data_in(a_data_8_4_to_8_5),
  .b_data_in(b_data_7_5_to_8_5),
  .c_data(c_data_8_5),
  .a_data_out(a_data_8_5_to_8_6),
  .b_data_out(b_data_8_5_to_9_5),
  .a_addr(a_addr_8_5_NC),
  .b_addr(b_addr_8_5_NC),
  .c_addr(c_addr_8_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 8_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_6_to_8_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_6_to_9_6;
  wire [`AWIDTH-1:0] a_addr_8_6_NC;
  wire [`AWIDTH-1:0] b_addr_8_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_6),
  .a_data(a_data_8_6_NC),
  .b_data(b_data_8_6_NC),
  .a_data_in(a_data_8_5_to_8_6),
  .b_data_in(b_data_7_6_to_8_6),
  .c_data(c_data_8_6),
  .a_data_out(a_data_8_6_to_8_7),
  .b_data_out(b_data_8_6_to_9_6),
  .a_addr(a_addr_8_6_NC),
  .b_addr(b_addr_8_6_NC),
  .c_addr(c_addr_8_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 8_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_7_to_8_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_7_to_9_7;
  wire [`AWIDTH-1:0] a_addr_8_7_NC;
  wire [`AWIDTH-1:0] b_addr_8_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_7),
  .a_data(a_data_8_7_NC),
  .b_data(b_data_8_7_NC),
  .a_data_in(a_data_8_6_to_8_7),
  .b_data_in(b_data_7_7_to_8_7),
  .c_data(c_data_8_7),
  .a_data_out(a_data_8_7_to_8_8),
  .b_data_out(b_data_8_7_to_9_7),
  .a_addr(a_addr_8_7_NC),
  .b_addr(b_addr_8_7_NC),
  .c_addr(c_addr_8_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 8_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_8_to_8_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_8_to_9_8;
  wire [`AWIDTH-1:0] a_addr_8_8_NC;
  wire [`AWIDTH-1:0] b_addr_8_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_8),
  .a_data(a_data_8_8_NC),
  .b_data(b_data_8_8_NC),
  .a_data_in(a_data_8_7_to_8_8),
  .b_data_in(b_data_7_8_to_8_8),
  .c_data(c_data_8_8),
  .a_data_out(a_data_8_8_to_8_9),
  .b_data_out(b_data_8_8_to_9_8),
  .a_addr(a_addr_8_8_NC),
  .b_addr(b_addr_8_8_NC),
  .c_addr(c_addr_8_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 8_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_9_to_8_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_9_to_9_9;
  wire [`AWIDTH-1:0] a_addr_8_9_NC;
  wire [`AWIDTH-1:0] b_addr_8_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_9),
  .a_data(a_data_8_9_NC),
  .b_data(b_data_8_9_NC),
  .a_data_in(a_data_8_8_to_8_9),
  .b_data_in(b_data_7_9_to_8_9),
  .c_data(c_data_8_9),
  .a_data_out(a_data_8_9_to_8_10),
  .b_data_out(b_data_8_9_to_9_9),
  .a_addr(a_addr_8_9_NC),
  .b_addr(b_addr_8_9_NC),
  .c_addr(c_addr_8_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 8_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_10_to_8_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_10_to_9_10;
  wire [`AWIDTH-1:0] a_addr_8_10_NC;
  wire [`AWIDTH-1:0] b_addr_8_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_10),
  .a_data(a_data_8_10_NC),
  .b_data(b_data_8_10_NC),
  .a_data_in(a_data_8_9_to_8_10),
  .b_data_in(b_data_7_10_to_8_10),
  .c_data(c_data_8_10),
  .a_data_out(a_data_8_10_to_8_11),
  .b_data_out(b_data_8_10_to_9_10),
  .a_addr(a_addr_8_10_NC),
  .b_addr(b_addr_8_10_NC),
  .c_addr(c_addr_8_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 8_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_11_to_8_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_11_to_9_11;
  wire [`AWIDTH-1:0] a_addr_8_11_NC;
  wire [`AWIDTH-1:0] b_addr_8_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_11),
  .a_data(a_data_8_11_NC),
  .b_data(b_data_8_11_NC),
  .a_data_in(a_data_8_10_to_8_11),
  .b_data_in(b_data_7_11_to_8_11),
  .c_data(c_data_8_11),
  .a_data_out(a_data_8_11_to_8_12),
  .b_data_out(b_data_8_11_to_9_11),
  .a_addr(a_addr_8_11_NC),
  .b_addr(b_addr_8_11_NC),
  .c_addr(c_addr_8_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 8_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_12_to_8_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_12_to_9_12;
  wire [`AWIDTH-1:0] a_addr_8_12_NC;
  wire [`AWIDTH-1:0] b_addr_8_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_12),
  .a_data(a_data_8_12_NC),
  .b_data(b_data_8_12_NC),
  .a_data_in(a_data_8_11_to_8_12),
  .b_data_in(b_data_7_12_to_8_12),
  .c_data(c_data_8_12),
  .a_data_out(a_data_8_12_to_8_13),
  .b_data_out(b_data_8_12_to_9_12),
  .a_addr(a_addr_8_12_NC),
  .b_addr(b_addr_8_12_NC),
  .c_addr(c_addr_8_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 8_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_13_to_8_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_13_to_9_13;
  wire [`AWIDTH-1:0] a_addr_8_13_NC;
  wire [`AWIDTH-1:0] b_addr_8_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_13),
  .a_data(a_data_8_13_NC),
  .b_data(b_data_8_13_NC),
  .a_data_in(a_data_8_12_to_8_13),
  .b_data_in(b_data_7_13_to_8_13),
  .c_data(c_data_8_13),
  .a_data_out(a_data_8_13_to_8_14),
  .b_data_out(b_data_8_13_to_9_13),
  .a_addr(a_addr_8_13_NC),
  .b_addr(b_addr_8_13_NC),
  .c_addr(c_addr_8_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 8_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_14_to_8_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_14_to_9_14;
  wire [`AWIDTH-1:0] a_addr_8_14_NC;
  wire [`AWIDTH-1:0] b_addr_8_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_14),
  .a_data(a_data_8_14_NC),
  .b_data(b_data_8_14_NC),
  .a_data_in(a_data_8_13_to_8_14),
  .b_data_in(b_data_7_14_to_8_14),
  .c_data(c_data_8_14),
  .a_data_out(a_data_8_14_to_8_15),
  .b_data_out(b_data_8_14_to_9_14),
  .a_addr(a_addr_8_14_NC),
  .b_addr(b_addr_8_14_NC),
  .c_addr(c_addr_8_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 8_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_15_to_8_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_15_to_9_15;
  wire [`AWIDTH-1:0] a_addr_8_15_NC;
  wire [`AWIDTH-1:0] b_addr_8_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_8_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_8_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_8_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_8_15),
  .a_data(a_data_8_15_NC),
  .b_data(b_data_8_15_NC),
  .a_data_in(a_data_8_14_to_8_15),
  .b_data_in(b_data_7_15_to_8_15),
  .c_data(c_data_8_15),
  .a_data_out(a_data_8_15_to_8_16),
  .b_data_out(b_data_8_15_to_9_15),
  .a_addr(a_addr_8_15_NC),
  .b_addr(b_addr_8_15_NC),
  .c_addr(c_addr_8_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd8),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 9_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_0_to_9_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_0_to_10_0;
  wire [`AWIDTH-1:0] b_addr_9_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_9_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_0),
  .a_data(a_data_9_0),
  .b_data(b_data_9_0_NC),
  .a_data_in(a_data_in_9_0_NC),
  .b_data_in(b_data_8_0_to_9_0),
  .c_data(c_data_9_0),
  .a_data_out(a_data_9_0_to_9_1),
  .b_data_out(b_data_9_0_to_10_0),
  .a_addr(a_addr_9_0),
  .b_addr(b_addr_9_0_NC),
  .c_addr(c_addr_9_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 9_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_1_to_9_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_1_to_10_1;
  wire [`AWIDTH-1:0] a_addr_9_1_NC;
  wire [`AWIDTH-1:0] b_addr_9_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_1),
  .a_data(a_data_9_1_NC),
  .b_data(b_data_9_1_NC),
  .a_data_in(a_data_9_0_to_9_1),
  .b_data_in(b_data_8_1_to_9_1),
  .c_data(c_data_9_1),
  .a_data_out(a_data_9_1_to_9_2),
  .b_data_out(b_data_9_1_to_10_1),
  .a_addr(a_addr_9_1_NC),
  .b_addr(b_addr_9_1_NC),
  .c_addr(c_addr_9_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 9_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_2_to_9_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_2_to_10_2;
  wire [`AWIDTH-1:0] a_addr_9_2_NC;
  wire [`AWIDTH-1:0] b_addr_9_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_2),
  .a_data(a_data_9_2_NC),
  .b_data(b_data_9_2_NC),
  .a_data_in(a_data_9_1_to_9_2),
  .b_data_in(b_data_8_2_to_9_2),
  .c_data(c_data_9_2),
  .a_data_out(a_data_9_2_to_9_3),
  .b_data_out(b_data_9_2_to_10_2),
  .a_addr(a_addr_9_2_NC),
  .b_addr(b_addr_9_2_NC),
  .c_addr(c_addr_9_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 9_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_3_to_9_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_3_to_10_3;
  wire [`AWIDTH-1:0] a_addr_9_3_NC;
  wire [`AWIDTH-1:0] b_addr_9_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_3),
  .a_data(a_data_9_3_NC),
  .b_data(b_data_9_3_NC),
  .a_data_in(a_data_9_2_to_9_3),
  .b_data_in(b_data_8_3_to_9_3),
  .c_data(c_data_9_3),
  .a_data_out(a_data_9_3_to_9_4),
  .b_data_out(b_data_9_3_to_10_3),
  .a_addr(a_addr_9_3_NC),
  .b_addr(b_addr_9_3_NC),
  .c_addr(c_addr_9_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 9_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_4_to_9_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_4_to_10_4;
  wire [`AWIDTH-1:0] a_addr_9_4_NC;
  wire [`AWIDTH-1:0] b_addr_9_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_4),
  .a_data(a_data_9_4_NC),
  .b_data(b_data_9_4_NC),
  .a_data_in(a_data_9_3_to_9_4),
  .b_data_in(b_data_8_4_to_9_4),
  .c_data(c_data_9_4),
  .a_data_out(a_data_9_4_to_9_5),
  .b_data_out(b_data_9_4_to_10_4),
  .a_addr(a_addr_9_4_NC),
  .b_addr(b_addr_9_4_NC),
  .c_addr(c_addr_9_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 9_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_5_to_9_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_5_to_10_5;
  wire [`AWIDTH-1:0] a_addr_9_5_NC;
  wire [`AWIDTH-1:0] b_addr_9_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_5),
  .a_data(a_data_9_5_NC),
  .b_data(b_data_9_5_NC),
  .a_data_in(a_data_9_4_to_9_5),
  .b_data_in(b_data_8_5_to_9_5),
  .c_data(c_data_9_5),
  .a_data_out(a_data_9_5_to_9_6),
  .b_data_out(b_data_9_5_to_10_5),
  .a_addr(a_addr_9_5_NC),
  .b_addr(b_addr_9_5_NC),
  .c_addr(c_addr_9_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 9_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_6_to_9_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_6_to_10_6;
  wire [`AWIDTH-1:0] a_addr_9_6_NC;
  wire [`AWIDTH-1:0] b_addr_9_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_6),
  .a_data(a_data_9_6_NC),
  .b_data(b_data_9_6_NC),
  .a_data_in(a_data_9_5_to_9_6),
  .b_data_in(b_data_8_6_to_9_6),
  .c_data(c_data_9_6),
  .a_data_out(a_data_9_6_to_9_7),
  .b_data_out(b_data_9_6_to_10_6),
  .a_addr(a_addr_9_6_NC),
  .b_addr(b_addr_9_6_NC),
  .c_addr(c_addr_9_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 9_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_7_to_9_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_7_to_10_7;
  wire [`AWIDTH-1:0] a_addr_9_7_NC;
  wire [`AWIDTH-1:0] b_addr_9_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_7),
  .a_data(a_data_9_7_NC),
  .b_data(b_data_9_7_NC),
  .a_data_in(a_data_9_6_to_9_7),
  .b_data_in(b_data_8_7_to_9_7),
  .c_data(c_data_9_7),
  .a_data_out(a_data_9_7_to_9_8),
  .b_data_out(b_data_9_7_to_10_7),
  .a_addr(a_addr_9_7_NC),
  .b_addr(b_addr_9_7_NC),
  .c_addr(c_addr_9_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 9_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_8_to_9_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_8_to_10_8;
  wire [`AWIDTH-1:0] a_addr_9_8_NC;
  wire [`AWIDTH-1:0] b_addr_9_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_8),
  .a_data(a_data_9_8_NC),
  .b_data(b_data_9_8_NC),
  .a_data_in(a_data_9_7_to_9_8),
  .b_data_in(b_data_8_8_to_9_8),
  .c_data(c_data_9_8),
  .a_data_out(a_data_9_8_to_9_9),
  .b_data_out(b_data_9_8_to_10_8),
  .a_addr(a_addr_9_8_NC),
  .b_addr(b_addr_9_8_NC),
  .c_addr(c_addr_9_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 9_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_9_to_9_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_9_to_10_9;
  wire [`AWIDTH-1:0] a_addr_9_9_NC;
  wire [`AWIDTH-1:0] b_addr_9_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_9),
  .a_data(a_data_9_9_NC),
  .b_data(b_data_9_9_NC),
  .a_data_in(a_data_9_8_to_9_9),
  .b_data_in(b_data_8_9_to_9_9),
  .c_data(c_data_9_9),
  .a_data_out(a_data_9_9_to_9_10),
  .b_data_out(b_data_9_9_to_10_9),
  .a_addr(a_addr_9_9_NC),
  .b_addr(b_addr_9_9_NC),
  .c_addr(c_addr_9_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 9_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_10_to_9_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_10_to_10_10;
  wire [`AWIDTH-1:0] a_addr_9_10_NC;
  wire [`AWIDTH-1:0] b_addr_9_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_10),
  .a_data(a_data_9_10_NC),
  .b_data(b_data_9_10_NC),
  .a_data_in(a_data_9_9_to_9_10),
  .b_data_in(b_data_8_10_to_9_10),
  .c_data(c_data_9_10),
  .a_data_out(a_data_9_10_to_9_11),
  .b_data_out(b_data_9_10_to_10_10),
  .a_addr(a_addr_9_10_NC),
  .b_addr(b_addr_9_10_NC),
  .c_addr(c_addr_9_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 9_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_11_to_9_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_11_to_10_11;
  wire [`AWIDTH-1:0] a_addr_9_11_NC;
  wire [`AWIDTH-1:0] b_addr_9_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_11),
  .a_data(a_data_9_11_NC),
  .b_data(b_data_9_11_NC),
  .a_data_in(a_data_9_10_to_9_11),
  .b_data_in(b_data_8_11_to_9_11),
  .c_data(c_data_9_11),
  .a_data_out(a_data_9_11_to_9_12),
  .b_data_out(b_data_9_11_to_10_11),
  .a_addr(a_addr_9_11_NC),
  .b_addr(b_addr_9_11_NC),
  .c_addr(c_addr_9_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 9_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_12_to_9_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_12_to_10_12;
  wire [`AWIDTH-1:0] a_addr_9_12_NC;
  wire [`AWIDTH-1:0] b_addr_9_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_12),
  .a_data(a_data_9_12_NC),
  .b_data(b_data_9_12_NC),
  .a_data_in(a_data_9_11_to_9_12),
  .b_data_in(b_data_8_12_to_9_12),
  .c_data(c_data_9_12),
  .a_data_out(a_data_9_12_to_9_13),
  .b_data_out(b_data_9_12_to_10_12),
  .a_addr(a_addr_9_12_NC),
  .b_addr(b_addr_9_12_NC),
  .c_addr(c_addr_9_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 9_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_13_to_9_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_13_to_10_13;
  wire [`AWIDTH-1:0] a_addr_9_13_NC;
  wire [`AWIDTH-1:0] b_addr_9_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_13),
  .a_data(a_data_9_13_NC),
  .b_data(b_data_9_13_NC),
  .a_data_in(a_data_9_12_to_9_13),
  .b_data_in(b_data_8_13_to_9_13),
  .c_data(c_data_9_13),
  .a_data_out(a_data_9_13_to_9_14),
  .b_data_out(b_data_9_13_to_10_13),
  .a_addr(a_addr_9_13_NC),
  .b_addr(b_addr_9_13_NC),
  .c_addr(c_addr_9_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 9_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_14_to_9_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_14_to_10_14;
  wire [`AWIDTH-1:0] a_addr_9_14_NC;
  wire [`AWIDTH-1:0] b_addr_9_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_14),
  .a_data(a_data_9_14_NC),
  .b_data(b_data_9_14_NC),
  .a_data_in(a_data_9_13_to_9_14),
  .b_data_in(b_data_8_14_to_9_14),
  .c_data(c_data_9_14),
  .a_data_out(a_data_9_14_to_9_15),
  .b_data_out(b_data_9_14_to_10_14),
  .a_addr(a_addr_9_14_NC),
  .b_addr(b_addr_9_14_NC),
  .c_addr(c_addr_9_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 9_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_15_to_9_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_15_to_10_15;
  wire [`AWIDTH-1:0] a_addr_9_15_NC;
  wire [`AWIDTH-1:0] b_addr_9_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_9_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_9_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_9_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_9_15),
  .a_data(a_data_9_15_NC),
  .b_data(b_data_9_15_NC),
  .a_data_in(a_data_9_14_to_9_15),
  .b_data_in(b_data_8_15_to_9_15),
  .c_data(c_data_9_15),
  .a_data_out(a_data_9_15_to_9_16),
  .b_data_out(b_data_9_15_to_10_15),
  .a_addr(a_addr_9_15_NC),
  .b_addr(b_addr_9_15_NC),
  .c_addr(c_addr_9_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd9),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 10_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_0_to_10_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_0_to_11_0;
  wire [`AWIDTH-1:0] b_addr_10_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_10_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_0),
  .a_data(a_data_10_0),
  .b_data(b_data_10_0_NC),
  .a_data_in(a_data_in_10_0_NC),
  .b_data_in(b_data_9_0_to_10_0),
  .c_data(c_data_10_0),
  .a_data_out(a_data_10_0_to_10_1),
  .b_data_out(b_data_10_0_to_11_0),
  .a_addr(a_addr_10_0),
  .b_addr(b_addr_10_0_NC),
  .c_addr(c_addr_10_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 10_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_1_to_10_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_1_to_11_1;
  wire [`AWIDTH-1:0] a_addr_10_1_NC;
  wire [`AWIDTH-1:0] b_addr_10_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_1),
  .a_data(a_data_10_1_NC),
  .b_data(b_data_10_1_NC),
  .a_data_in(a_data_10_0_to_10_1),
  .b_data_in(b_data_9_1_to_10_1),
  .c_data(c_data_10_1),
  .a_data_out(a_data_10_1_to_10_2),
  .b_data_out(b_data_10_1_to_11_1),
  .a_addr(a_addr_10_1_NC),
  .b_addr(b_addr_10_1_NC),
  .c_addr(c_addr_10_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 10_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_2_to_10_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_2_to_11_2;
  wire [`AWIDTH-1:0] a_addr_10_2_NC;
  wire [`AWIDTH-1:0] b_addr_10_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_2),
  .a_data(a_data_10_2_NC),
  .b_data(b_data_10_2_NC),
  .a_data_in(a_data_10_1_to_10_2),
  .b_data_in(b_data_9_2_to_10_2),
  .c_data(c_data_10_2),
  .a_data_out(a_data_10_2_to_10_3),
  .b_data_out(b_data_10_2_to_11_2),
  .a_addr(a_addr_10_2_NC),
  .b_addr(b_addr_10_2_NC),
  .c_addr(c_addr_10_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 10_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_3_to_10_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_3_to_11_3;
  wire [`AWIDTH-1:0] a_addr_10_3_NC;
  wire [`AWIDTH-1:0] b_addr_10_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_3),
  .a_data(a_data_10_3_NC),
  .b_data(b_data_10_3_NC),
  .a_data_in(a_data_10_2_to_10_3),
  .b_data_in(b_data_9_3_to_10_3),
  .c_data(c_data_10_3),
  .a_data_out(a_data_10_3_to_10_4),
  .b_data_out(b_data_10_3_to_11_3),
  .a_addr(a_addr_10_3_NC),
  .b_addr(b_addr_10_3_NC),
  .c_addr(c_addr_10_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 10_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_4_to_10_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_4_to_11_4;
  wire [`AWIDTH-1:0] a_addr_10_4_NC;
  wire [`AWIDTH-1:0] b_addr_10_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_4),
  .a_data(a_data_10_4_NC),
  .b_data(b_data_10_4_NC),
  .a_data_in(a_data_10_3_to_10_4),
  .b_data_in(b_data_9_4_to_10_4),
  .c_data(c_data_10_4),
  .a_data_out(a_data_10_4_to_10_5),
  .b_data_out(b_data_10_4_to_11_4),
  .a_addr(a_addr_10_4_NC),
  .b_addr(b_addr_10_4_NC),
  .c_addr(c_addr_10_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 10_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_5_to_10_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_5_to_11_5;
  wire [`AWIDTH-1:0] a_addr_10_5_NC;
  wire [`AWIDTH-1:0] b_addr_10_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_5),
  .a_data(a_data_10_5_NC),
  .b_data(b_data_10_5_NC),
  .a_data_in(a_data_10_4_to_10_5),
  .b_data_in(b_data_9_5_to_10_5),
  .c_data(c_data_10_5),
  .a_data_out(a_data_10_5_to_10_6),
  .b_data_out(b_data_10_5_to_11_5),
  .a_addr(a_addr_10_5_NC),
  .b_addr(b_addr_10_5_NC),
  .c_addr(c_addr_10_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 10_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_6_to_10_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_6_to_11_6;
  wire [`AWIDTH-1:0] a_addr_10_6_NC;
  wire [`AWIDTH-1:0] b_addr_10_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_6),
  .a_data(a_data_10_6_NC),
  .b_data(b_data_10_6_NC),
  .a_data_in(a_data_10_5_to_10_6),
  .b_data_in(b_data_9_6_to_10_6),
  .c_data(c_data_10_6),
  .a_data_out(a_data_10_6_to_10_7),
  .b_data_out(b_data_10_6_to_11_6),
  .a_addr(a_addr_10_6_NC),
  .b_addr(b_addr_10_6_NC),
  .c_addr(c_addr_10_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 10_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_7_to_10_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_7_to_11_7;
  wire [`AWIDTH-1:0] a_addr_10_7_NC;
  wire [`AWIDTH-1:0] b_addr_10_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_7),
  .a_data(a_data_10_7_NC),
  .b_data(b_data_10_7_NC),
  .a_data_in(a_data_10_6_to_10_7),
  .b_data_in(b_data_9_7_to_10_7),
  .c_data(c_data_10_7),
  .a_data_out(a_data_10_7_to_10_8),
  .b_data_out(b_data_10_7_to_11_7),
  .a_addr(a_addr_10_7_NC),
  .b_addr(b_addr_10_7_NC),
  .c_addr(c_addr_10_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 10_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_8_to_10_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_8_to_11_8;
  wire [`AWIDTH-1:0] a_addr_10_8_NC;
  wire [`AWIDTH-1:0] b_addr_10_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_8),
  .a_data(a_data_10_8_NC),
  .b_data(b_data_10_8_NC),
  .a_data_in(a_data_10_7_to_10_8),
  .b_data_in(b_data_9_8_to_10_8),
  .c_data(c_data_10_8),
  .a_data_out(a_data_10_8_to_10_9),
  .b_data_out(b_data_10_8_to_11_8),
  .a_addr(a_addr_10_8_NC),
  .b_addr(b_addr_10_8_NC),
  .c_addr(c_addr_10_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 10_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_9_to_10_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_9_to_11_9;
  wire [`AWIDTH-1:0] a_addr_10_9_NC;
  wire [`AWIDTH-1:0] b_addr_10_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_9),
  .a_data(a_data_10_9_NC),
  .b_data(b_data_10_9_NC),
  .a_data_in(a_data_10_8_to_10_9),
  .b_data_in(b_data_9_9_to_10_9),
  .c_data(c_data_10_9),
  .a_data_out(a_data_10_9_to_10_10),
  .b_data_out(b_data_10_9_to_11_9),
  .a_addr(a_addr_10_9_NC),
  .b_addr(b_addr_10_9_NC),
  .c_addr(c_addr_10_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 10_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_10_to_10_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_10_to_11_10;
  wire [`AWIDTH-1:0] a_addr_10_10_NC;
  wire [`AWIDTH-1:0] b_addr_10_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_10),
  .a_data(a_data_10_10_NC),
  .b_data(b_data_10_10_NC),
  .a_data_in(a_data_10_9_to_10_10),
  .b_data_in(b_data_9_10_to_10_10),
  .c_data(c_data_10_10),
  .a_data_out(a_data_10_10_to_10_11),
  .b_data_out(b_data_10_10_to_11_10),
  .a_addr(a_addr_10_10_NC),
  .b_addr(b_addr_10_10_NC),
  .c_addr(c_addr_10_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 10_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_11_to_10_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_11_to_11_11;
  wire [`AWIDTH-1:0] a_addr_10_11_NC;
  wire [`AWIDTH-1:0] b_addr_10_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_11),
  .a_data(a_data_10_11_NC),
  .b_data(b_data_10_11_NC),
  .a_data_in(a_data_10_10_to_10_11),
  .b_data_in(b_data_9_11_to_10_11),
  .c_data(c_data_10_11),
  .a_data_out(a_data_10_11_to_10_12),
  .b_data_out(b_data_10_11_to_11_11),
  .a_addr(a_addr_10_11_NC),
  .b_addr(b_addr_10_11_NC),
  .c_addr(c_addr_10_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 10_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_12_to_10_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_12_to_11_12;
  wire [`AWIDTH-1:0] a_addr_10_12_NC;
  wire [`AWIDTH-1:0] b_addr_10_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_12),
  .a_data(a_data_10_12_NC),
  .b_data(b_data_10_12_NC),
  .a_data_in(a_data_10_11_to_10_12),
  .b_data_in(b_data_9_12_to_10_12),
  .c_data(c_data_10_12),
  .a_data_out(a_data_10_12_to_10_13),
  .b_data_out(b_data_10_12_to_11_12),
  .a_addr(a_addr_10_12_NC),
  .b_addr(b_addr_10_12_NC),
  .c_addr(c_addr_10_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 10_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_13_to_10_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_13_to_11_13;
  wire [`AWIDTH-1:0] a_addr_10_13_NC;
  wire [`AWIDTH-1:0] b_addr_10_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_13),
  .a_data(a_data_10_13_NC),
  .b_data(b_data_10_13_NC),
  .a_data_in(a_data_10_12_to_10_13),
  .b_data_in(b_data_9_13_to_10_13),
  .c_data(c_data_10_13),
  .a_data_out(a_data_10_13_to_10_14),
  .b_data_out(b_data_10_13_to_11_13),
  .a_addr(a_addr_10_13_NC),
  .b_addr(b_addr_10_13_NC),
  .c_addr(c_addr_10_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 10_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_14_to_10_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_14_to_11_14;
  wire [`AWIDTH-1:0] a_addr_10_14_NC;
  wire [`AWIDTH-1:0] b_addr_10_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_14),
  .a_data(a_data_10_14_NC),
  .b_data(b_data_10_14_NC),
  .a_data_in(a_data_10_13_to_10_14),
  .b_data_in(b_data_9_14_to_10_14),
  .c_data(c_data_10_14),
  .a_data_out(a_data_10_14_to_10_15),
  .b_data_out(b_data_10_14_to_11_14),
  .a_addr(a_addr_10_14_NC),
  .b_addr(b_addr_10_14_NC),
  .c_addr(c_addr_10_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 10_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_15_to_10_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_15_to_11_15;
  wire [`AWIDTH-1:0] a_addr_10_15_NC;
  wire [`AWIDTH-1:0] b_addr_10_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_10_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_10_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_10_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_10_15),
  .a_data(a_data_10_15_NC),
  .b_data(b_data_10_15_NC),
  .a_data_in(a_data_10_14_to_10_15),
  .b_data_in(b_data_9_15_to_10_15),
  .c_data(c_data_10_15),
  .a_data_out(a_data_10_15_to_10_16),
  .b_data_out(b_data_10_15_to_11_15),
  .a_addr(a_addr_10_15_NC),
  .b_addr(b_addr_10_15_NC),
  .c_addr(c_addr_10_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd10),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 11_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_0_to_11_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_0_to_12_0;
  wire [`AWIDTH-1:0] b_addr_11_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_11_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_0),
  .a_data(a_data_11_0),
  .b_data(b_data_11_0_NC),
  .a_data_in(a_data_in_11_0_NC),
  .b_data_in(b_data_10_0_to_11_0),
  .c_data(c_data_11_0),
  .a_data_out(a_data_11_0_to_11_1),
  .b_data_out(b_data_11_0_to_12_0),
  .a_addr(a_addr_11_0),
  .b_addr(b_addr_11_0_NC),
  .c_addr(c_addr_11_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 11_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_1_to_11_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_1_to_12_1;
  wire [`AWIDTH-1:0] a_addr_11_1_NC;
  wire [`AWIDTH-1:0] b_addr_11_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_1),
  .a_data(a_data_11_1_NC),
  .b_data(b_data_11_1_NC),
  .a_data_in(a_data_11_0_to_11_1),
  .b_data_in(b_data_10_1_to_11_1),
  .c_data(c_data_11_1),
  .a_data_out(a_data_11_1_to_11_2),
  .b_data_out(b_data_11_1_to_12_1),
  .a_addr(a_addr_11_1_NC),
  .b_addr(b_addr_11_1_NC),
  .c_addr(c_addr_11_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 11_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_2_to_11_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_2_to_12_2;
  wire [`AWIDTH-1:0] a_addr_11_2_NC;
  wire [`AWIDTH-1:0] b_addr_11_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_2),
  .a_data(a_data_11_2_NC),
  .b_data(b_data_11_2_NC),
  .a_data_in(a_data_11_1_to_11_2),
  .b_data_in(b_data_10_2_to_11_2),
  .c_data(c_data_11_2),
  .a_data_out(a_data_11_2_to_11_3),
  .b_data_out(b_data_11_2_to_12_2),
  .a_addr(a_addr_11_2_NC),
  .b_addr(b_addr_11_2_NC),
  .c_addr(c_addr_11_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 11_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_3_to_11_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_3_to_12_3;
  wire [`AWIDTH-1:0] a_addr_11_3_NC;
  wire [`AWIDTH-1:0] b_addr_11_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_3),
  .a_data(a_data_11_3_NC),
  .b_data(b_data_11_3_NC),
  .a_data_in(a_data_11_2_to_11_3),
  .b_data_in(b_data_10_3_to_11_3),
  .c_data(c_data_11_3),
  .a_data_out(a_data_11_3_to_11_4),
  .b_data_out(b_data_11_3_to_12_3),
  .a_addr(a_addr_11_3_NC),
  .b_addr(b_addr_11_3_NC),
  .c_addr(c_addr_11_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 11_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_4_to_11_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_4_to_12_4;
  wire [`AWIDTH-1:0] a_addr_11_4_NC;
  wire [`AWIDTH-1:0] b_addr_11_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_4),
  .a_data(a_data_11_4_NC),
  .b_data(b_data_11_4_NC),
  .a_data_in(a_data_11_3_to_11_4),
  .b_data_in(b_data_10_4_to_11_4),
  .c_data(c_data_11_4),
  .a_data_out(a_data_11_4_to_11_5),
  .b_data_out(b_data_11_4_to_12_4),
  .a_addr(a_addr_11_4_NC),
  .b_addr(b_addr_11_4_NC),
  .c_addr(c_addr_11_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 11_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_5_to_11_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_5_to_12_5;
  wire [`AWIDTH-1:0] a_addr_11_5_NC;
  wire [`AWIDTH-1:0] b_addr_11_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_5),
  .a_data(a_data_11_5_NC),
  .b_data(b_data_11_5_NC),
  .a_data_in(a_data_11_4_to_11_5),
  .b_data_in(b_data_10_5_to_11_5),
  .c_data(c_data_11_5),
  .a_data_out(a_data_11_5_to_11_6),
  .b_data_out(b_data_11_5_to_12_5),
  .a_addr(a_addr_11_5_NC),
  .b_addr(b_addr_11_5_NC),
  .c_addr(c_addr_11_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 11_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_6_to_11_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_6_to_12_6;
  wire [`AWIDTH-1:0] a_addr_11_6_NC;
  wire [`AWIDTH-1:0] b_addr_11_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_6),
  .a_data(a_data_11_6_NC),
  .b_data(b_data_11_6_NC),
  .a_data_in(a_data_11_5_to_11_6),
  .b_data_in(b_data_10_6_to_11_6),
  .c_data(c_data_11_6),
  .a_data_out(a_data_11_6_to_11_7),
  .b_data_out(b_data_11_6_to_12_6),
  .a_addr(a_addr_11_6_NC),
  .b_addr(b_addr_11_6_NC),
  .c_addr(c_addr_11_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 11_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_7_to_11_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_7_to_12_7;
  wire [`AWIDTH-1:0] a_addr_11_7_NC;
  wire [`AWIDTH-1:0] b_addr_11_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_7),
  .a_data(a_data_11_7_NC),
  .b_data(b_data_11_7_NC),
  .a_data_in(a_data_11_6_to_11_7),
  .b_data_in(b_data_10_7_to_11_7),
  .c_data(c_data_11_7),
  .a_data_out(a_data_11_7_to_11_8),
  .b_data_out(b_data_11_7_to_12_7),
  .a_addr(a_addr_11_7_NC),
  .b_addr(b_addr_11_7_NC),
  .c_addr(c_addr_11_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 11_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_8_to_11_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_8_to_12_8;
  wire [`AWIDTH-1:0] a_addr_11_8_NC;
  wire [`AWIDTH-1:0] b_addr_11_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_8),
  .a_data(a_data_11_8_NC),
  .b_data(b_data_11_8_NC),
  .a_data_in(a_data_11_7_to_11_8),
  .b_data_in(b_data_10_8_to_11_8),
  .c_data(c_data_11_8),
  .a_data_out(a_data_11_8_to_11_9),
  .b_data_out(b_data_11_8_to_12_8),
  .a_addr(a_addr_11_8_NC),
  .b_addr(b_addr_11_8_NC),
  .c_addr(c_addr_11_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 11_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_9_to_11_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_9_to_12_9;
  wire [`AWIDTH-1:0] a_addr_11_9_NC;
  wire [`AWIDTH-1:0] b_addr_11_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_9),
  .a_data(a_data_11_9_NC),
  .b_data(b_data_11_9_NC),
  .a_data_in(a_data_11_8_to_11_9),
  .b_data_in(b_data_10_9_to_11_9),
  .c_data(c_data_11_9),
  .a_data_out(a_data_11_9_to_11_10),
  .b_data_out(b_data_11_9_to_12_9),
  .a_addr(a_addr_11_9_NC),
  .b_addr(b_addr_11_9_NC),
  .c_addr(c_addr_11_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 11_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_10_to_11_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_10_to_12_10;
  wire [`AWIDTH-1:0] a_addr_11_10_NC;
  wire [`AWIDTH-1:0] b_addr_11_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_10),
  .a_data(a_data_11_10_NC),
  .b_data(b_data_11_10_NC),
  .a_data_in(a_data_11_9_to_11_10),
  .b_data_in(b_data_10_10_to_11_10),
  .c_data(c_data_11_10),
  .a_data_out(a_data_11_10_to_11_11),
  .b_data_out(b_data_11_10_to_12_10),
  .a_addr(a_addr_11_10_NC),
  .b_addr(b_addr_11_10_NC),
  .c_addr(c_addr_11_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 11_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_11_to_11_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_11_to_12_11;
  wire [`AWIDTH-1:0] a_addr_11_11_NC;
  wire [`AWIDTH-1:0] b_addr_11_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_11),
  .a_data(a_data_11_11_NC),
  .b_data(b_data_11_11_NC),
  .a_data_in(a_data_11_10_to_11_11),
  .b_data_in(b_data_10_11_to_11_11),
  .c_data(c_data_11_11),
  .a_data_out(a_data_11_11_to_11_12),
  .b_data_out(b_data_11_11_to_12_11),
  .a_addr(a_addr_11_11_NC),
  .b_addr(b_addr_11_11_NC),
  .c_addr(c_addr_11_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 11_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_12_to_11_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_12_to_12_12;
  wire [`AWIDTH-1:0] a_addr_11_12_NC;
  wire [`AWIDTH-1:0] b_addr_11_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_12),
  .a_data(a_data_11_12_NC),
  .b_data(b_data_11_12_NC),
  .a_data_in(a_data_11_11_to_11_12),
  .b_data_in(b_data_10_12_to_11_12),
  .c_data(c_data_11_12),
  .a_data_out(a_data_11_12_to_11_13),
  .b_data_out(b_data_11_12_to_12_12),
  .a_addr(a_addr_11_12_NC),
  .b_addr(b_addr_11_12_NC),
  .c_addr(c_addr_11_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 11_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_13_to_11_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_13_to_12_13;
  wire [`AWIDTH-1:0] a_addr_11_13_NC;
  wire [`AWIDTH-1:0] b_addr_11_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_13),
  .a_data(a_data_11_13_NC),
  .b_data(b_data_11_13_NC),
  .a_data_in(a_data_11_12_to_11_13),
  .b_data_in(b_data_10_13_to_11_13),
  .c_data(c_data_11_13),
  .a_data_out(a_data_11_13_to_11_14),
  .b_data_out(b_data_11_13_to_12_13),
  .a_addr(a_addr_11_13_NC),
  .b_addr(b_addr_11_13_NC),
  .c_addr(c_addr_11_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 11_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_14_to_11_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_14_to_12_14;
  wire [`AWIDTH-1:0] a_addr_11_14_NC;
  wire [`AWIDTH-1:0] b_addr_11_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_14),
  .a_data(a_data_11_14_NC),
  .b_data(b_data_11_14_NC),
  .a_data_in(a_data_11_13_to_11_14),
  .b_data_in(b_data_10_14_to_11_14),
  .c_data(c_data_11_14),
  .a_data_out(a_data_11_14_to_11_15),
  .b_data_out(b_data_11_14_to_12_14),
  .a_addr(a_addr_11_14_NC),
  .b_addr(b_addr_11_14_NC),
  .c_addr(c_addr_11_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 11_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_15_to_11_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_15_to_12_15;
  wire [`AWIDTH-1:0] a_addr_11_15_NC;
  wire [`AWIDTH-1:0] b_addr_11_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_11_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_11_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_11_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_11_15),
  .a_data(a_data_11_15_NC),
  .b_data(b_data_11_15_NC),
  .a_data_in(a_data_11_14_to_11_15),
  .b_data_in(b_data_10_15_to_11_15),
  .c_data(c_data_11_15),
  .a_data_out(a_data_11_15_to_11_16),
  .b_data_out(b_data_11_15_to_12_15),
  .a_addr(a_addr_11_15_NC),
  .b_addr(b_addr_11_15_NC),
  .c_addr(c_addr_11_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd11),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 12_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_0_to_12_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_0_to_13_0;
  wire [`AWIDTH-1:0] b_addr_12_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_12_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_0),
  .a_data(a_data_12_0),
  .b_data(b_data_12_0_NC),
  .a_data_in(a_data_in_12_0_NC),
  .b_data_in(b_data_11_0_to_12_0),
  .c_data(c_data_12_0),
  .a_data_out(a_data_12_0_to_12_1),
  .b_data_out(b_data_12_0_to_13_0),
  .a_addr(a_addr_12_0),
  .b_addr(b_addr_12_0_NC),
  .c_addr(c_addr_12_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 12_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_1_to_12_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_1_to_13_1;
  wire [`AWIDTH-1:0] a_addr_12_1_NC;
  wire [`AWIDTH-1:0] b_addr_12_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_1),
  .a_data(a_data_12_1_NC),
  .b_data(b_data_12_1_NC),
  .a_data_in(a_data_12_0_to_12_1),
  .b_data_in(b_data_11_1_to_12_1),
  .c_data(c_data_12_1),
  .a_data_out(a_data_12_1_to_12_2),
  .b_data_out(b_data_12_1_to_13_1),
  .a_addr(a_addr_12_1_NC),
  .b_addr(b_addr_12_1_NC),
  .c_addr(c_addr_12_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 12_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_2_to_12_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_2_to_13_2;
  wire [`AWIDTH-1:0] a_addr_12_2_NC;
  wire [`AWIDTH-1:0] b_addr_12_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_2),
  .a_data(a_data_12_2_NC),
  .b_data(b_data_12_2_NC),
  .a_data_in(a_data_12_1_to_12_2),
  .b_data_in(b_data_11_2_to_12_2),
  .c_data(c_data_12_2),
  .a_data_out(a_data_12_2_to_12_3),
  .b_data_out(b_data_12_2_to_13_2),
  .a_addr(a_addr_12_2_NC),
  .b_addr(b_addr_12_2_NC),
  .c_addr(c_addr_12_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 12_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_3_to_12_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_3_to_13_3;
  wire [`AWIDTH-1:0] a_addr_12_3_NC;
  wire [`AWIDTH-1:0] b_addr_12_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_3),
  .a_data(a_data_12_3_NC),
  .b_data(b_data_12_3_NC),
  .a_data_in(a_data_12_2_to_12_3),
  .b_data_in(b_data_11_3_to_12_3),
  .c_data(c_data_12_3),
  .a_data_out(a_data_12_3_to_12_4),
  .b_data_out(b_data_12_3_to_13_3),
  .a_addr(a_addr_12_3_NC),
  .b_addr(b_addr_12_3_NC),
  .c_addr(c_addr_12_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 12_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_4_to_12_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_4_to_13_4;
  wire [`AWIDTH-1:0] a_addr_12_4_NC;
  wire [`AWIDTH-1:0] b_addr_12_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_4),
  .a_data(a_data_12_4_NC),
  .b_data(b_data_12_4_NC),
  .a_data_in(a_data_12_3_to_12_4),
  .b_data_in(b_data_11_4_to_12_4),
  .c_data(c_data_12_4),
  .a_data_out(a_data_12_4_to_12_5),
  .b_data_out(b_data_12_4_to_13_4),
  .a_addr(a_addr_12_4_NC),
  .b_addr(b_addr_12_4_NC),
  .c_addr(c_addr_12_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 12_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_5_to_12_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_5_to_13_5;
  wire [`AWIDTH-1:0] a_addr_12_5_NC;
  wire [`AWIDTH-1:0] b_addr_12_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_5),
  .a_data(a_data_12_5_NC),
  .b_data(b_data_12_5_NC),
  .a_data_in(a_data_12_4_to_12_5),
  .b_data_in(b_data_11_5_to_12_5),
  .c_data(c_data_12_5),
  .a_data_out(a_data_12_5_to_12_6),
  .b_data_out(b_data_12_5_to_13_5),
  .a_addr(a_addr_12_5_NC),
  .b_addr(b_addr_12_5_NC),
  .c_addr(c_addr_12_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 12_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_6_to_12_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_6_to_13_6;
  wire [`AWIDTH-1:0] a_addr_12_6_NC;
  wire [`AWIDTH-1:0] b_addr_12_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_6),
  .a_data(a_data_12_6_NC),
  .b_data(b_data_12_6_NC),
  .a_data_in(a_data_12_5_to_12_6),
  .b_data_in(b_data_11_6_to_12_6),
  .c_data(c_data_12_6),
  .a_data_out(a_data_12_6_to_12_7),
  .b_data_out(b_data_12_6_to_13_6),
  .a_addr(a_addr_12_6_NC),
  .b_addr(b_addr_12_6_NC),
  .c_addr(c_addr_12_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 12_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_7_to_12_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_7_to_13_7;
  wire [`AWIDTH-1:0] a_addr_12_7_NC;
  wire [`AWIDTH-1:0] b_addr_12_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_7),
  .a_data(a_data_12_7_NC),
  .b_data(b_data_12_7_NC),
  .a_data_in(a_data_12_6_to_12_7),
  .b_data_in(b_data_11_7_to_12_7),
  .c_data(c_data_12_7),
  .a_data_out(a_data_12_7_to_12_8),
  .b_data_out(b_data_12_7_to_13_7),
  .a_addr(a_addr_12_7_NC),
  .b_addr(b_addr_12_7_NC),
  .c_addr(c_addr_12_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 12_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_8_to_12_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_8_to_13_8;
  wire [`AWIDTH-1:0] a_addr_12_8_NC;
  wire [`AWIDTH-1:0] b_addr_12_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_8),
  .a_data(a_data_12_8_NC),
  .b_data(b_data_12_8_NC),
  .a_data_in(a_data_12_7_to_12_8),
  .b_data_in(b_data_11_8_to_12_8),
  .c_data(c_data_12_8),
  .a_data_out(a_data_12_8_to_12_9),
  .b_data_out(b_data_12_8_to_13_8),
  .a_addr(a_addr_12_8_NC),
  .b_addr(b_addr_12_8_NC),
  .c_addr(c_addr_12_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 12_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_9_to_12_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_9_to_13_9;
  wire [`AWIDTH-1:0] a_addr_12_9_NC;
  wire [`AWIDTH-1:0] b_addr_12_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_9),
  .a_data(a_data_12_9_NC),
  .b_data(b_data_12_9_NC),
  .a_data_in(a_data_12_8_to_12_9),
  .b_data_in(b_data_11_9_to_12_9),
  .c_data(c_data_12_9),
  .a_data_out(a_data_12_9_to_12_10),
  .b_data_out(b_data_12_9_to_13_9),
  .a_addr(a_addr_12_9_NC),
  .b_addr(b_addr_12_9_NC),
  .c_addr(c_addr_12_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 12_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_10_to_12_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_10_to_13_10;
  wire [`AWIDTH-1:0] a_addr_12_10_NC;
  wire [`AWIDTH-1:0] b_addr_12_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_10),
  .a_data(a_data_12_10_NC),
  .b_data(b_data_12_10_NC),
  .a_data_in(a_data_12_9_to_12_10),
  .b_data_in(b_data_11_10_to_12_10),
  .c_data(c_data_12_10),
  .a_data_out(a_data_12_10_to_12_11),
  .b_data_out(b_data_12_10_to_13_10),
  .a_addr(a_addr_12_10_NC),
  .b_addr(b_addr_12_10_NC),
  .c_addr(c_addr_12_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 12_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_11_to_12_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_11_to_13_11;
  wire [`AWIDTH-1:0] a_addr_12_11_NC;
  wire [`AWIDTH-1:0] b_addr_12_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_11),
  .a_data(a_data_12_11_NC),
  .b_data(b_data_12_11_NC),
  .a_data_in(a_data_12_10_to_12_11),
  .b_data_in(b_data_11_11_to_12_11),
  .c_data(c_data_12_11),
  .a_data_out(a_data_12_11_to_12_12),
  .b_data_out(b_data_12_11_to_13_11),
  .a_addr(a_addr_12_11_NC),
  .b_addr(b_addr_12_11_NC),
  .c_addr(c_addr_12_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 12_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_12_to_12_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_12_to_13_12;
  wire [`AWIDTH-1:0] a_addr_12_12_NC;
  wire [`AWIDTH-1:0] b_addr_12_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_12),
  .a_data(a_data_12_12_NC),
  .b_data(b_data_12_12_NC),
  .a_data_in(a_data_12_11_to_12_12),
  .b_data_in(b_data_11_12_to_12_12),
  .c_data(c_data_12_12),
  .a_data_out(a_data_12_12_to_12_13),
  .b_data_out(b_data_12_12_to_13_12),
  .a_addr(a_addr_12_12_NC),
  .b_addr(b_addr_12_12_NC),
  .c_addr(c_addr_12_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 12_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_13_to_12_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_13_to_13_13;
  wire [`AWIDTH-1:0] a_addr_12_13_NC;
  wire [`AWIDTH-1:0] b_addr_12_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_13),
  .a_data(a_data_12_13_NC),
  .b_data(b_data_12_13_NC),
  .a_data_in(a_data_12_12_to_12_13),
  .b_data_in(b_data_11_13_to_12_13),
  .c_data(c_data_12_13),
  .a_data_out(a_data_12_13_to_12_14),
  .b_data_out(b_data_12_13_to_13_13),
  .a_addr(a_addr_12_13_NC),
  .b_addr(b_addr_12_13_NC),
  .c_addr(c_addr_12_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 12_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_14_to_12_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_14_to_13_14;
  wire [`AWIDTH-1:0] a_addr_12_14_NC;
  wire [`AWIDTH-1:0] b_addr_12_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_14),
  .a_data(a_data_12_14_NC),
  .b_data(b_data_12_14_NC),
  .a_data_in(a_data_12_13_to_12_14),
  .b_data_in(b_data_11_14_to_12_14),
  .c_data(c_data_12_14),
  .a_data_out(a_data_12_14_to_12_15),
  .b_data_out(b_data_12_14_to_13_14),
  .a_addr(a_addr_12_14_NC),
  .b_addr(b_addr_12_14_NC),
  .c_addr(c_addr_12_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 12_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_15_to_12_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_15_to_13_15;
  wire [`AWIDTH-1:0] a_addr_12_15_NC;
  wire [`AWIDTH-1:0] b_addr_12_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_12_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_12_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_12_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_12_15),
  .a_data(a_data_12_15_NC),
  .b_data(b_data_12_15_NC),
  .a_data_in(a_data_12_14_to_12_15),
  .b_data_in(b_data_11_15_to_12_15),
  .c_data(c_data_12_15),
  .a_data_out(a_data_12_15_to_12_16),
  .b_data_out(b_data_12_15_to_13_15),
  .a_addr(a_addr_12_15_NC),
  .b_addr(b_addr_12_15_NC),
  .c_addr(c_addr_12_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd12),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 13_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_0_to_13_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_0_to_14_0;
  wire [`AWIDTH-1:0] b_addr_13_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_13_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_0),
  .a_data(a_data_13_0),
  .b_data(b_data_13_0_NC),
  .a_data_in(a_data_in_13_0_NC),
  .b_data_in(b_data_12_0_to_13_0),
  .c_data(c_data_13_0),
  .a_data_out(a_data_13_0_to_13_1),
  .b_data_out(b_data_13_0_to_14_0),
  .a_addr(a_addr_13_0),
  .b_addr(b_addr_13_0_NC),
  .c_addr(c_addr_13_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 13_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_1_to_13_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_1_to_14_1;
  wire [`AWIDTH-1:0] a_addr_13_1_NC;
  wire [`AWIDTH-1:0] b_addr_13_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_1),
  .a_data(a_data_13_1_NC),
  .b_data(b_data_13_1_NC),
  .a_data_in(a_data_13_0_to_13_1),
  .b_data_in(b_data_12_1_to_13_1),
  .c_data(c_data_13_1),
  .a_data_out(a_data_13_1_to_13_2),
  .b_data_out(b_data_13_1_to_14_1),
  .a_addr(a_addr_13_1_NC),
  .b_addr(b_addr_13_1_NC),
  .c_addr(c_addr_13_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 13_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_2_to_13_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_2_to_14_2;
  wire [`AWIDTH-1:0] a_addr_13_2_NC;
  wire [`AWIDTH-1:0] b_addr_13_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_2),
  .a_data(a_data_13_2_NC),
  .b_data(b_data_13_2_NC),
  .a_data_in(a_data_13_1_to_13_2),
  .b_data_in(b_data_12_2_to_13_2),
  .c_data(c_data_13_2),
  .a_data_out(a_data_13_2_to_13_3),
  .b_data_out(b_data_13_2_to_14_2),
  .a_addr(a_addr_13_2_NC),
  .b_addr(b_addr_13_2_NC),
  .c_addr(c_addr_13_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 13_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_3_to_13_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_3_to_14_3;
  wire [`AWIDTH-1:0] a_addr_13_3_NC;
  wire [`AWIDTH-1:0] b_addr_13_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_3),
  .a_data(a_data_13_3_NC),
  .b_data(b_data_13_3_NC),
  .a_data_in(a_data_13_2_to_13_3),
  .b_data_in(b_data_12_3_to_13_3),
  .c_data(c_data_13_3),
  .a_data_out(a_data_13_3_to_13_4),
  .b_data_out(b_data_13_3_to_14_3),
  .a_addr(a_addr_13_3_NC),
  .b_addr(b_addr_13_3_NC),
  .c_addr(c_addr_13_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 13_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_4_to_13_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_4_to_14_4;
  wire [`AWIDTH-1:0] a_addr_13_4_NC;
  wire [`AWIDTH-1:0] b_addr_13_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_4),
  .a_data(a_data_13_4_NC),
  .b_data(b_data_13_4_NC),
  .a_data_in(a_data_13_3_to_13_4),
  .b_data_in(b_data_12_4_to_13_4),
  .c_data(c_data_13_4),
  .a_data_out(a_data_13_4_to_13_5),
  .b_data_out(b_data_13_4_to_14_4),
  .a_addr(a_addr_13_4_NC),
  .b_addr(b_addr_13_4_NC),
  .c_addr(c_addr_13_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 13_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_5_to_13_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_5_to_14_5;
  wire [`AWIDTH-1:0] a_addr_13_5_NC;
  wire [`AWIDTH-1:0] b_addr_13_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_5),
  .a_data(a_data_13_5_NC),
  .b_data(b_data_13_5_NC),
  .a_data_in(a_data_13_4_to_13_5),
  .b_data_in(b_data_12_5_to_13_5),
  .c_data(c_data_13_5),
  .a_data_out(a_data_13_5_to_13_6),
  .b_data_out(b_data_13_5_to_14_5),
  .a_addr(a_addr_13_5_NC),
  .b_addr(b_addr_13_5_NC),
  .c_addr(c_addr_13_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 13_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_6_to_13_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_6_to_14_6;
  wire [`AWIDTH-1:0] a_addr_13_6_NC;
  wire [`AWIDTH-1:0] b_addr_13_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_6),
  .a_data(a_data_13_6_NC),
  .b_data(b_data_13_6_NC),
  .a_data_in(a_data_13_5_to_13_6),
  .b_data_in(b_data_12_6_to_13_6),
  .c_data(c_data_13_6),
  .a_data_out(a_data_13_6_to_13_7),
  .b_data_out(b_data_13_6_to_14_6),
  .a_addr(a_addr_13_6_NC),
  .b_addr(b_addr_13_6_NC),
  .c_addr(c_addr_13_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 13_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_7_to_13_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_7_to_14_7;
  wire [`AWIDTH-1:0] a_addr_13_7_NC;
  wire [`AWIDTH-1:0] b_addr_13_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_7),
  .a_data(a_data_13_7_NC),
  .b_data(b_data_13_7_NC),
  .a_data_in(a_data_13_6_to_13_7),
  .b_data_in(b_data_12_7_to_13_7),
  .c_data(c_data_13_7),
  .a_data_out(a_data_13_7_to_13_8),
  .b_data_out(b_data_13_7_to_14_7),
  .a_addr(a_addr_13_7_NC),
  .b_addr(b_addr_13_7_NC),
  .c_addr(c_addr_13_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 13_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_8_to_13_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_8_to_14_8;
  wire [`AWIDTH-1:0] a_addr_13_8_NC;
  wire [`AWIDTH-1:0] b_addr_13_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_8),
  .a_data(a_data_13_8_NC),
  .b_data(b_data_13_8_NC),
  .a_data_in(a_data_13_7_to_13_8),
  .b_data_in(b_data_12_8_to_13_8),
  .c_data(c_data_13_8),
  .a_data_out(a_data_13_8_to_13_9),
  .b_data_out(b_data_13_8_to_14_8),
  .a_addr(a_addr_13_8_NC),
  .b_addr(b_addr_13_8_NC),
  .c_addr(c_addr_13_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 13_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_9_to_13_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_9_to_14_9;
  wire [`AWIDTH-1:0] a_addr_13_9_NC;
  wire [`AWIDTH-1:0] b_addr_13_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_9),
  .a_data(a_data_13_9_NC),
  .b_data(b_data_13_9_NC),
  .a_data_in(a_data_13_8_to_13_9),
  .b_data_in(b_data_12_9_to_13_9),
  .c_data(c_data_13_9),
  .a_data_out(a_data_13_9_to_13_10),
  .b_data_out(b_data_13_9_to_14_9),
  .a_addr(a_addr_13_9_NC),
  .b_addr(b_addr_13_9_NC),
  .c_addr(c_addr_13_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 13_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_10_to_13_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_10_to_14_10;
  wire [`AWIDTH-1:0] a_addr_13_10_NC;
  wire [`AWIDTH-1:0] b_addr_13_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_10),
  .a_data(a_data_13_10_NC),
  .b_data(b_data_13_10_NC),
  .a_data_in(a_data_13_9_to_13_10),
  .b_data_in(b_data_12_10_to_13_10),
  .c_data(c_data_13_10),
  .a_data_out(a_data_13_10_to_13_11),
  .b_data_out(b_data_13_10_to_14_10),
  .a_addr(a_addr_13_10_NC),
  .b_addr(b_addr_13_10_NC),
  .c_addr(c_addr_13_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 13_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_11_to_13_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_11_to_14_11;
  wire [`AWIDTH-1:0] a_addr_13_11_NC;
  wire [`AWIDTH-1:0] b_addr_13_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_11),
  .a_data(a_data_13_11_NC),
  .b_data(b_data_13_11_NC),
  .a_data_in(a_data_13_10_to_13_11),
  .b_data_in(b_data_12_11_to_13_11),
  .c_data(c_data_13_11),
  .a_data_out(a_data_13_11_to_13_12),
  .b_data_out(b_data_13_11_to_14_11),
  .a_addr(a_addr_13_11_NC),
  .b_addr(b_addr_13_11_NC),
  .c_addr(c_addr_13_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 13_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_12_to_13_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_12_to_14_12;
  wire [`AWIDTH-1:0] a_addr_13_12_NC;
  wire [`AWIDTH-1:0] b_addr_13_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_12),
  .a_data(a_data_13_12_NC),
  .b_data(b_data_13_12_NC),
  .a_data_in(a_data_13_11_to_13_12),
  .b_data_in(b_data_12_12_to_13_12),
  .c_data(c_data_13_12),
  .a_data_out(a_data_13_12_to_13_13),
  .b_data_out(b_data_13_12_to_14_12),
  .a_addr(a_addr_13_12_NC),
  .b_addr(b_addr_13_12_NC),
  .c_addr(c_addr_13_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 13_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_13_to_13_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_13_to_14_13;
  wire [`AWIDTH-1:0] a_addr_13_13_NC;
  wire [`AWIDTH-1:0] b_addr_13_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_13),
  .a_data(a_data_13_13_NC),
  .b_data(b_data_13_13_NC),
  .a_data_in(a_data_13_12_to_13_13),
  .b_data_in(b_data_12_13_to_13_13),
  .c_data(c_data_13_13),
  .a_data_out(a_data_13_13_to_13_14),
  .b_data_out(b_data_13_13_to_14_13),
  .a_addr(a_addr_13_13_NC),
  .b_addr(b_addr_13_13_NC),
  .c_addr(c_addr_13_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 13_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_14_to_13_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_14_to_14_14;
  wire [`AWIDTH-1:0] a_addr_13_14_NC;
  wire [`AWIDTH-1:0] b_addr_13_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_14),
  .a_data(a_data_13_14_NC),
  .b_data(b_data_13_14_NC),
  .a_data_in(a_data_13_13_to_13_14),
  .b_data_in(b_data_12_14_to_13_14),
  .c_data(c_data_13_14),
  .a_data_out(a_data_13_14_to_13_15),
  .b_data_out(b_data_13_14_to_14_14),
  .a_addr(a_addr_13_14_NC),
  .b_addr(b_addr_13_14_NC),
  .c_addr(c_addr_13_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 13_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_15_to_13_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_15_to_14_15;
  wire [`AWIDTH-1:0] a_addr_13_15_NC;
  wire [`AWIDTH-1:0] b_addr_13_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_13_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_13_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_13_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_13_15),
  .a_data(a_data_13_15_NC),
  .b_data(b_data_13_15_NC),
  .a_data_in(a_data_13_14_to_13_15),
  .b_data_in(b_data_12_15_to_13_15),
  .c_data(c_data_13_15),
  .a_data_out(a_data_13_15_to_13_16),
  .b_data_out(b_data_13_15_to_14_15),
  .a_addr(a_addr_13_15_NC),
  .b_addr(b_addr_13_15_NC),
  .c_addr(c_addr_13_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd13),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 14_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_0_to_14_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_0_to_15_0;
  wire [`AWIDTH-1:0] b_addr_14_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_14_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_0),
  .a_data(a_data_14_0),
  .b_data(b_data_14_0_NC),
  .a_data_in(a_data_in_14_0_NC),
  .b_data_in(b_data_13_0_to_14_0),
  .c_data(c_data_14_0),
  .a_data_out(a_data_14_0_to_14_1),
  .b_data_out(b_data_14_0_to_15_0),
  .a_addr(a_addr_14_0),
  .b_addr(b_addr_14_0_NC),
  .c_addr(c_addr_14_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 14_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_1_to_14_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_1_to_15_1;
  wire [`AWIDTH-1:0] a_addr_14_1_NC;
  wire [`AWIDTH-1:0] b_addr_14_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_1),
  .a_data(a_data_14_1_NC),
  .b_data(b_data_14_1_NC),
  .a_data_in(a_data_14_0_to_14_1),
  .b_data_in(b_data_13_1_to_14_1),
  .c_data(c_data_14_1),
  .a_data_out(a_data_14_1_to_14_2),
  .b_data_out(b_data_14_1_to_15_1),
  .a_addr(a_addr_14_1_NC),
  .b_addr(b_addr_14_1_NC),
  .c_addr(c_addr_14_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 14_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_2_to_14_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_2_to_15_2;
  wire [`AWIDTH-1:0] a_addr_14_2_NC;
  wire [`AWIDTH-1:0] b_addr_14_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_2),
  .a_data(a_data_14_2_NC),
  .b_data(b_data_14_2_NC),
  .a_data_in(a_data_14_1_to_14_2),
  .b_data_in(b_data_13_2_to_14_2),
  .c_data(c_data_14_2),
  .a_data_out(a_data_14_2_to_14_3),
  .b_data_out(b_data_14_2_to_15_2),
  .a_addr(a_addr_14_2_NC),
  .b_addr(b_addr_14_2_NC),
  .c_addr(c_addr_14_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 14_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_3_to_14_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_3_to_15_3;
  wire [`AWIDTH-1:0] a_addr_14_3_NC;
  wire [`AWIDTH-1:0] b_addr_14_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_3),
  .a_data(a_data_14_3_NC),
  .b_data(b_data_14_3_NC),
  .a_data_in(a_data_14_2_to_14_3),
  .b_data_in(b_data_13_3_to_14_3),
  .c_data(c_data_14_3),
  .a_data_out(a_data_14_3_to_14_4),
  .b_data_out(b_data_14_3_to_15_3),
  .a_addr(a_addr_14_3_NC),
  .b_addr(b_addr_14_3_NC),
  .c_addr(c_addr_14_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 14_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_4_to_14_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_4_to_15_4;
  wire [`AWIDTH-1:0] a_addr_14_4_NC;
  wire [`AWIDTH-1:0] b_addr_14_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_4),
  .a_data(a_data_14_4_NC),
  .b_data(b_data_14_4_NC),
  .a_data_in(a_data_14_3_to_14_4),
  .b_data_in(b_data_13_4_to_14_4),
  .c_data(c_data_14_4),
  .a_data_out(a_data_14_4_to_14_5),
  .b_data_out(b_data_14_4_to_15_4),
  .a_addr(a_addr_14_4_NC),
  .b_addr(b_addr_14_4_NC),
  .c_addr(c_addr_14_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 14_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_5_to_14_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_5_to_15_5;
  wire [`AWIDTH-1:0] a_addr_14_5_NC;
  wire [`AWIDTH-1:0] b_addr_14_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_5),
  .a_data(a_data_14_5_NC),
  .b_data(b_data_14_5_NC),
  .a_data_in(a_data_14_4_to_14_5),
  .b_data_in(b_data_13_5_to_14_5),
  .c_data(c_data_14_5),
  .a_data_out(a_data_14_5_to_14_6),
  .b_data_out(b_data_14_5_to_15_5),
  .a_addr(a_addr_14_5_NC),
  .b_addr(b_addr_14_5_NC),
  .c_addr(c_addr_14_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 14_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_6_to_14_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_6_to_15_6;
  wire [`AWIDTH-1:0] a_addr_14_6_NC;
  wire [`AWIDTH-1:0] b_addr_14_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_6),
  .a_data(a_data_14_6_NC),
  .b_data(b_data_14_6_NC),
  .a_data_in(a_data_14_5_to_14_6),
  .b_data_in(b_data_13_6_to_14_6),
  .c_data(c_data_14_6),
  .a_data_out(a_data_14_6_to_14_7),
  .b_data_out(b_data_14_6_to_15_6),
  .a_addr(a_addr_14_6_NC),
  .b_addr(b_addr_14_6_NC),
  .c_addr(c_addr_14_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 14_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_7_to_14_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_7_to_15_7;
  wire [`AWIDTH-1:0] a_addr_14_7_NC;
  wire [`AWIDTH-1:0] b_addr_14_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_7),
  .a_data(a_data_14_7_NC),
  .b_data(b_data_14_7_NC),
  .a_data_in(a_data_14_6_to_14_7),
  .b_data_in(b_data_13_7_to_14_7),
  .c_data(c_data_14_7),
  .a_data_out(a_data_14_7_to_14_8),
  .b_data_out(b_data_14_7_to_15_7),
  .a_addr(a_addr_14_7_NC),
  .b_addr(b_addr_14_7_NC),
  .c_addr(c_addr_14_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 14_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_8_to_14_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_8_to_15_8;
  wire [`AWIDTH-1:0] a_addr_14_8_NC;
  wire [`AWIDTH-1:0] b_addr_14_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_8),
  .a_data(a_data_14_8_NC),
  .b_data(b_data_14_8_NC),
  .a_data_in(a_data_14_7_to_14_8),
  .b_data_in(b_data_13_8_to_14_8),
  .c_data(c_data_14_8),
  .a_data_out(a_data_14_8_to_14_9),
  .b_data_out(b_data_14_8_to_15_8),
  .a_addr(a_addr_14_8_NC),
  .b_addr(b_addr_14_8_NC),
  .c_addr(c_addr_14_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 14_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_9_to_14_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_9_to_15_9;
  wire [`AWIDTH-1:0] a_addr_14_9_NC;
  wire [`AWIDTH-1:0] b_addr_14_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_9),
  .a_data(a_data_14_9_NC),
  .b_data(b_data_14_9_NC),
  .a_data_in(a_data_14_8_to_14_9),
  .b_data_in(b_data_13_9_to_14_9),
  .c_data(c_data_14_9),
  .a_data_out(a_data_14_9_to_14_10),
  .b_data_out(b_data_14_9_to_15_9),
  .a_addr(a_addr_14_9_NC),
  .b_addr(b_addr_14_9_NC),
  .c_addr(c_addr_14_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 14_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_10_to_14_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_10_to_15_10;
  wire [`AWIDTH-1:0] a_addr_14_10_NC;
  wire [`AWIDTH-1:0] b_addr_14_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_10),
  .a_data(a_data_14_10_NC),
  .b_data(b_data_14_10_NC),
  .a_data_in(a_data_14_9_to_14_10),
  .b_data_in(b_data_13_10_to_14_10),
  .c_data(c_data_14_10),
  .a_data_out(a_data_14_10_to_14_11),
  .b_data_out(b_data_14_10_to_15_10),
  .a_addr(a_addr_14_10_NC),
  .b_addr(b_addr_14_10_NC),
  .c_addr(c_addr_14_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 14_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_11_to_14_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_11_to_15_11;
  wire [`AWIDTH-1:0] a_addr_14_11_NC;
  wire [`AWIDTH-1:0] b_addr_14_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_11),
  .a_data(a_data_14_11_NC),
  .b_data(b_data_14_11_NC),
  .a_data_in(a_data_14_10_to_14_11),
  .b_data_in(b_data_13_11_to_14_11),
  .c_data(c_data_14_11),
  .a_data_out(a_data_14_11_to_14_12),
  .b_data_out(b_data_14_11_to_15_11),
  .a_addr(a_addr_14_11_NC),
  .b_addr(b_addr_14_11_NC),
  .c_addr(c_addr_14_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 14_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_12_to_14_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_12_to_15_12;
  wire [`AWIDTH-1:0] a_addr_14_12_NC;
  wire [`AWIDTH-1:0] b_addr_14_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_12),
  .a_data(a_data_14_12_NC),
  .b_data(b_data_14_12_NC),
  .a_data_in(a_data_14_11_to_14_12),
  .b_data_in(b_data_13_12_to_14_12),
  .c_data(c_data_14_12),
  .a_data_out(a_data_14_12_to_14_13),
  .b_data_out(b_data_14_12_to_15_12),
  .a_addr(a_addr_14_12_NC),
  .b_addr(b_addr_14_12_NC),
  .c_addr(c_addr_14_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 14_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_13_to_14_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_13_to_15_13;
  wire [`AWIDTH-1:0] a_addr_14_13_NC;
  wire [`AWIDTH-1:0] b_addr_14_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_13),
  .a_data(a_data_14_13_NC),
  .b_data(b_data_14_13_NC),
  .a_data_in(a_data_14_12_to_14_13),
  .b_data_in(b_data_13_13_to_14_13),
  .c_data(c_data_14_13),
  .a_data_out(a_data_14_13_to_14_14),
  .b_data_out(b_data_14_13_to_15_13),
  .a_addr(a_addr_14_13_NC),
  .b_addr(b_addr_14_13_NC),
  .c_addr(c_addr_14_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 14_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_14_to_14_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_14_to_15_14;
  wire [`AWIDTH-1:0] a_addr_14_14_NC;
  wire [`AWIDTH-1:0] b_addr_14_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_14),
  .a_data(a_data_14_14_NC),
  .b_data(b_data_14_14_NC),
  .a_data_in(a_data_14_13_to_14_14),
  .b_data_in(b_data_13_14_to_14_14),
  .c_data(c_data_14_14),
  .a_data_out(a_data_14_14_to_14_15),
  .b_data_out(b_data_14_14_to_15_14),
  .a_addr(a_addr_14_14_NC),
  .b_addr(b_addr_14_14_NC),
  .c_addr(c_addr_14_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 14_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_15_to_14_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_15_to_15_15;
  wire [`AWIDTH-1:0] a_addr_14_15_NC;
  wire [`AWIDTH-1:0] b_addr_14_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_14_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_14_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_14_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_14_15),
  .a_data(a_data_14_15_NC),
  .b_data(b_data_14_15_NC),
  .a_data_in(a_data_14_14_to_14_15),
  .b_data_in(b_data_13_15_to_14_15),
  .c_data(c_data_14_15),
  .a_data_out(a_data_14_15_to_14_16),
  .b_data_out(b_data_14_15_to_15_15),
  .a_addr(a_addr_14_15_NC),
  .b_addr(b_addr_14_15_NC),
  .c_addr(c_addr_14_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd14),
  .b_loc(8'd15)
);

  /////////////////////////////////////////////////
  // Matmul 15_0
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_0_to_15_1;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_0_to_16_0;
  wire [`AWIDTH-1:0] b_addr_15_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_0_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in_15_0_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_0(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_0),
  .a_data(a_data_15_0),
  .b_data(b_data_15_0_NC),
  .a_data_in(a_data_in_15_0_NC),
  .b_data_in(b_data_14_0_to_15_0),
  .c_data(c_data_15_0),
  .a_data_out(a_data_15_0_to_15_1),
  .b_data_out(b_data_15_0_to_16_0),
  .a_addr(a_addr_15_0),
  .b_addr(b_addr_15_0_NC),
  .c_addr(c_addr_15_0),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd0)
);

  /////////////////////////////////////////////////
  // Matmul 15_1
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_1_to_15_2;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_1_to_16_1;
  wire [`AWIDTH-1:0] a_addr_15_1_NC;
  wire [`AWIDTH-1:0] b_addr_15_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_1_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_1_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_1(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_1),
  .a_data(a_data_15_1_NC),
  .b_data(b_data_15_1_NC),
  .a_data_in(a_data_15_0_to_15_1),
  .b_data_in(b_data_14_1_to_15_1),
  .c_data(c_data_15_1),
  .a_data_out(a_data_15_1_to_15_2),
  .b_data_out(b_data_15_1_to_16_1),
  .a_addr(a_addr_15_1_NC),
  .b_addr(b_addr_15_1_NC),
  .c_addr(c_addr_15_1),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd1)
);

  /////////////////////////////////////////////////
  // Matmul 15_2
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_2_to_15_3;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_2_to_16_2;
  wire [`AWIDTH-1:0] a_addr_15_2_NC;
  wire [`AWIDTH-1:0] b_addr_15_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_2_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_2_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_2(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_2),
  .a_data(a_data_15_2_NC),
  .b_data(b_data_15_2_NC),
  .a_data_in(a_data_15_1_to_15_2),
  .b_data_in(b_data_14_2_to_15_2),
  .c_data(c_data_15_2),
  .a_data_out(a_data_15_2_to_15_3),
  .b_data_out(b_data_15_2_to_16_2),
  .a_addr(a_addr_15_2_NC),
  .b_addr(b_addr_15_2_NC),
  .c_addr(c_addr_15_2),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd2)
);

  /////////////////////////////////////////////////
  // Matmul 15_3
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_3_to_15_4;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_3_to_16_3;
  wire [`AWIDTH-1:0] a_addr_15_3_NC;
  wire [`AWIDTH-1:0] b_addr_15_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_3_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_3_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_3(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_3),
  .a_data(a_data_15_3_NC),
  .b_data(b_data_15_3_NC),
  .a_data_in(a_data_15_2_to_15_3),
  .b_data_in(b_data_14_3_to_15_3),
  .c_data(c_data_15_3),
  .a_data_out(a_data_15_3_to_15_4),
  .b_data_out(b_data_15_3_to_16_3),
  .a_addr(a_addr_15_3_NC),
  .b_addr(b_addr_15_3_NC),
  .c_addr(c_addr_15_3),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd3)
);

  /////////////////////////////////////////////////
  // Matmul 15_4
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_4_to_15_5;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_4_to_16_4;
  wire [`AWIDTH-1:0] a_addr_15_4_NC;
  wire [`AWIDTH-1:0] b_addr_15_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_4_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_4_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_4(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_4),
  .a_data(a_data_15_4_NC),
  .b_data(b_data_15_4_NC),
  .a_data_in(a_data_15_3_to_15_4),
  .b_data_in(b_data_14_4_to_15_4),
  .c_data(c_data_15_4),
  .a_data_out(a_data_15_4_to_15_5),
  .b_data_out(b_data_15_4_to_16_4),
  .a_addr(a_addr_15_4_NC),
  .b_addr(b_addr_15_4_NC),
  .c_addr(c_addr_15_4),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd4)
);

  /////////////////////////////////////////////////
  // Matmul 15_5
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_5_to_15_6;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_5_to_16_5;
  wire [`AWIDTH-1:0] a_addr_15_5_NC;
  wire [`AWIDTH-1:0] b_addr_15_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_5_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_5_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_5(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_5),
  .a_data(a_data_15_5_NC),
  .b_data(b_data_15_5_NC),
  .a_data_in(a_data_15_4_to_15_5),
  .b_data_in(b_data_14_5_to_15_5),
  .c_data(c_data_15_5),
  .a_data_out(a_data_15_5_to_15_6),
  .b_data_out(b_data_15_5_to_16_5),
  .a_addr(a_addr_15_5_NC),
  .b_addr(b_addr_15_5_NC),
  .c_addr(c_addr_15_5),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd5)
);

  /////////////////////////////////////////////////
  // Matmul 15_6
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_6_to_15_7;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_6_to_16_6;
  wire [`AWIDTH-1:0] a_addr_15_6_NC;
  wire [`AWIDTH-1:0] b_addr_15_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_6_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_6_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_6(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_6),
  .a_data(a_data_15_6_NC),
  .b_data(b_data_15_6_NC),
  .a_data_in(a_data_15_5_to_15_6),
  .b_data_in(b_data_14_6_to_15_6),
  .c_data(c_data_15_6),
  .a_data_out(a_data_15_6_to_15_7),
  .b_data_out(b_data_15_6_to_16_6),
  .a_addr(a_addr_15_6_NC),
  .b_addr(b_addr_15_6_NC),
  .c_addr(c_addr_15_6),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd6)
);

  /////////////////////////////////////////////////
  // Matmul 15_7
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_7_to_15_8;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_7_to_16_7;
  wire [`AWIDTH-1:0] a_addr_15_7_NC;
  wire [`AWIDTH-1:0] b_addr_15_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_7_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_7_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_7(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_7),
  .a_data(a_data_15_7_NC),
  .b_data(b_data_15_7_NC),
  .a_data_in(a_data_15_6_to_15_7),
  .b_data_in(b_data_14_7_to_15_7),
  .c_data(c_data_15_7),
  .a_data_out(a_data_15_7_to_15_8),
  .b_data_out(b_data_15_7_to_16_7),
  .a_addr(a_addr_15_7_NC),
  .b_addr(b_addr_15_7_NC),
  .c_addr(c_addr_15_7),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd7)
);

  /////////////////////////////////////////////////
  // Matmul 15_8
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_8_to_15_9;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_8_to_16_8;
  wire [`AWIDTH-1:0] a_addr_15_8_NC;
  wire [`AWIDTH-1:0] b_addr_15_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_8_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_8_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_8(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_8),
  .a_data(a_data_15_8_NC),
  .b_data(b_data_15_8_NC),
  .a_data_in(a_data_15_7_to_15_8),
  .b_data_in(b_data_14_8_to_15_8),
  .c_data(c_data_15_8),
  .a_data_out(a_data_15_8_to_15_9),
  .b_data_out(b_data_15_8_to_16_8),
  .a_addr(a_addr_15_8_NC),
  .b_addr(b_addr_15_8_NC),
  .c_addr(c_addr_15_8),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd8)
);

  /////////////////////////////////////////////////
  // Matmul 15_9
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_9_to_15_10;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_9_to_16_9;
  wire [`AWIDTH-1:0] a_addr_15_9_NC;
  wire [`AWIDTH-1:0] b_addr_15_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_9_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_9_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_9(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_9),
  .a_data(a_data_15_9_NC),
  .b_data(b_data_15_9_NC),
  .a_data_in(a_data_15_8_to_15_9),
  .b_data_in(b_data_14_9_to_15_9),
  .c_data(c_data_15_9),
  .a_data_out(a_data_15_9_to_15_10),
  .b_data_out(b_data_15_9_to_16_9),
  .a_addr(a_addr_15_9_NC),
  .b_addr(b_addr_15_9_NC),
  .c_addr(c_addr_15_9),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd9)
);

  /////////////////////////////////////////////////
  // Matmul 15_10
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_10_to_15_11;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_10_to_16_10;
  wire [`AWIDTH-1:0] a_addr_15_10_NC;
  wire [`AWIDTH-1:0] b_addr_15_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_10_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_10_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_10(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_10),
  .a_data(a_data_15_10_NC),
  .b_data(b_data_15_10_NC),
  .a_data_in(a_data_15_9_to_15_10),
  .b_data_in(b_data_14_10_to_15_10),
  .c_data(c_data_15_10),
  .a_data_out(a_data_15_10_to_15_11),
  .b_data_out(b_data_15_10_to_16_10),
  .a_addr(a_addr_15_10_NC),
  .b_addr(b_addr_15_10_NC),
  .c_addr(c_addr_15_10),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd10)
);

  /////////////////////////////////////////////////
  // Matmul 15_11
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_11_to_15_12;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_11_to_16_11;
  wire [`AWIDTH-1:0] a_addr_15_11_NC;
  wire [`AWIDTH-1:0] b_addr_15_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_11_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_11_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_11(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_11),
  .a_data(a_data_15_11_NC),
  .b_data(b_data_15_11_NC),
  .a_data_in(a_data_15_10_to_15_11),
  .b_data_in(b_data_14_11_to_15_11),
  .c_data(c_data_15_11),
  .a_data_out(a_data_15_11_to_15_12),
  .b_data_out(b_data_15_11_to_16_11),
  .a_addr(a_addr_15_11_NC),
  .b_addr(b_addr_15_11_NC),
  .c_addr(c_addr_15_11),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd11)
);

  /////////////////////////////////////////////////
  // Matmul 15_12
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_12_to_15_13;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_12_to_16_12;
  wire [`AWIDTH-1:0] a_addr_15_12_NC;
  wire [`AWIDTH-1:0] b_addr_15_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_12_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_12_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_12(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_12),
  .a_data(a_data_15_12_NC),
  .b_data(b_data_15_12_NC),
  .a_data_in(a_data_15_11_to_15_12),
  .b_data_in(b_data_14_12_to_15_12),
  .c_data(c_data_15_12),
  .a_data_out(a_data_15_12_to_15_13),
  .b_data_out(b_data_15_12_to_16_12),
  .a_addr(a_addr_15_12_NC),
  .b_addr(b_addr_15_12_NC),
  .c_addr(c_addr_15_12),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd12)
);

  /////////////////////////////////////////////////
  // Matmul 15_13
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_13_to_15_14;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_13_to_16_13;
  wire [`AWIDTH-1:0] a_addr_15_13_NC;
  wire [`AWIDTH-1:0] b_addr_15_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_13_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_13_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_13(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_13),
  .a_data(a_data_15_13_NC),
  .b_data(b_data_15_13_NC),
  .a_data_in(a_data_15_12_to_15_13),
  .b_data_in(b_data_14_13_to_15_13),
  .c_data(c_data_15_13),
  .a_data_out(a_data_15_13_to_15_14),
  .b_data_out(b_data_15_13_to_16_13),
  .a_addr(a_addr_15_13_NC),
  .b_addr(b_addr_15_13_NC),
  .c_addr(c_addr_15_13),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd13)
);

  /////////////////////////////////////////////////
  // Matmul 15_14
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_14_to_15_15;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_14_to_16_14;
  wire [`AWIDTH-1:0] a_addr_15_14_NC;
  wire [`AWIDTH-1:0] b_addr_15_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_14_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_14_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_14(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_14),
  .a_data(a_data_15_14_NC),
  .b_data(b_data_15_14_NC),
  .a_data_in(a_data_15_13_to_15_14),
  .b_data_in(b_data_14_14_to_15_14),
  .c_data(c_data_15_14),
  .a_data_out(a_data_15_14_to_15_15),
  .b_data_out(b_data_15_14_to_16_14),
  .a_addr(a_addr_15_14_NC),
  .b_addr(b_addr_15_14_NC),
  .c_addr(c_addr_15_14),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd14)
);

  /////////////////////////////////////////////////
  // Matmul 15_15
  /////////////////////////////////////////////////

  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_15_to_15_16;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_15_to_16_15;
  wire [`AWIDTH-1:0] a_addr_15_15_NC;
  wire [`AWIDTH-1:0] b_addr_15_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] a_data_15_15_NC;
  wire [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] b_data_15_15_NC;

matmul_4x4_systolic u_matmul_4x4_systolic_15_15(
  .clk(clk),
  .reset(reset),
  .start_mat_mul(start_mat_mul),
  .done_mat_mul(done_mat_mul_15_15),
  .a_data(a_data_15_15_NC),
  .b_data(b_data_15_15_NC),
  .a_data_in(a_data_15_14_to_15_15),
  .b_data_in(b_data_14_15_to_15_15),
  .c_data(c_data_15_15),
  .a_data_out(a_data_15_15_to_15_16),
  .b_data_out(b_data_15_15_to_16_15),
  .a_addr(a_addr_15_15_NC),
  .b_addr(b_addr_15_15_NC),
  .c_addr(c_addr_15_15),
  .final_mat_mul_size(8'd64),
  .a_loc(8'd15),
  .b_loc(8'd15)
);

endmodule

module ram (addr0, d0, we0, q0, clk);

input [`AWIDTH-1:0] addr0;
input [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] d0;
input we0;
output [`BB_MAT_MUL_SIZE*`DWIDTH-1:0] q0;
input clk;

single_port_ram u_single_port_ram(
  .data(d0),
  .we(we0),
  .addr(addr0),
  .clk(clk),
  .out(q0)
);
endmodule