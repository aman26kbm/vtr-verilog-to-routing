//////////////////////////////////////////////////////////////////////////////
//HLS generated design for 4-layered binary neural network 
//The dataflow is specific to the network
//The design uses 16-bit fixed point for activations, binary for weights 
//The dense layers are binary. Activation is relu.
//There is no memory, design uses registers to store activations and weights. 
//Generated from HLS using hls4ml
//The network used was https://github.com/fastmachinelearning/example-models/blob/master/keras/KERAS_3layer_binarydense_relu_max.json
//////////////////////////////////////////////////////////////////////////////

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

//////////////////////////////////////////////////////////////////////////////
// Abridged for VTR by: Aman Arora
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps 

module dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 (
        ap_clk,
        ap_rst,
        data_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [255:0] data_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
output  [15:0] ap_return_32;
output  [15:0] ap_return_33;
output  [15:0] ap_return_34;
output  [15:0] ap_return_35;
output  [15:0] ap_return_36;
output  [15:0] ap_return_37;
output  [15:0] ap_return_38;
output  [15:0] ap_return_39;
output  [15:0] ap_return_40;
output  [15:0] ap_return_41;
output  [15:0] ap_return_42;
output  [15:0] ap_return_43;
output  [15:0] ap_return_44;
output  [15:0] ap_return_45;
output  [15:0] ap_return_46;
output  [15:0] ap_return_47;
output  [15:0] ap_return_48;
output  [15:0] ap_return_49;
output  [15:0] ap_return_50;
output  [15:0] ap_return_51;
output  [15:0] ap_return_52;
output  [15:0] ap_return_53;
output  [15:0] ap_return_54;
output  [15:0] ap_return_55;
output  [15:0] ap_return_56;
output  [15:0] ap_return_57;
output  [15:0] ap_return_58;
output  [15:0] ap_return_59;
output  [15:0] ap_return_60;
output  [15:0] ap_return_61;
output  [15:0] ap_return_62;
output  [15:0] ap_return_63;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;
reg[15:0] ap_return_32;
reg[15:0] ap_return_33;
reg[15:0] ap_return_34;
reg[15:0] ap_return_35;
reg[15:0] ap_return_36;
reg[15:0] ap_return_37;
reg[15:0] ap_return_38;
reg[15:0] ap_return_39;
reg[15:0] ap_return_40;
reg[15:0] ap_return_41;
reg[15:0] ap_return_42;
reg[15:0] ap_return_43;
reg[15:0] ap_return_44;
reg[15:0] ap_return_45;
reg[15:0] ap_return_46;
reg[15:0] ap_return_47;
reg[15:0] ap_return_48;
reg[15:0] ap_return_49;
reg[15:0] ap_return_50;
reg[15:0] ap_return_51;
reg[15:0] ap_return_52;
reg[15:0] ap_return_53;
reg[15:0] ap_return_54;
reg[15:0] ap_return_55;
reg[15:0] ap_return_56;
reg[15:0] ap_return_57;
reg[15:0] ap_return_58;
reg[15:0] ap_return_59;
reg[15:0] ap_return_60;
reg[15:0] ap_return_61;
reg[15:0] ap_return_62;
reg[15:0] ap_return_63;

wire   [15:0] trunc_ln203_fu_88_p1;
reg   [15:0] trunc_ln203_reg_3431;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_pp0_stage0_11001;
wire   [15:0] tmp_2_fu_92_p4;
reg   [15:0] tmp_2_reg_3437;
reg   [15:0] tmp_3_reg_3443;
reg   [15:0] tmp_3_reg_3443_pp0_iter1_reg;
reg   [15:0] tmp_3_reg_3443_pp0_iter2_reg;
reg   [15:0] tmp_4_reg_3454;
reg   [15:0] tmp_4_reg_3454_pp0_iter1_reg;
reg   [15:0] tmp_4_reg_3454_pp0_iter2_reg;
reg   [15:0] tmp_4_reg_3454_pp0_iter3_reg;
reg   [15:0] tmp_4_reg_3454_pp0_iter4_reg;
reg   [15:0] mult_307_V_reg_3472;
reg   [15:0] mult_307_V_reg_3472_pp0_iter1_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter2_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter3_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter4_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter5_reg;
reg   [15:0] mult_320_V_reg_3500;
reg   [15:0] mult_320_V_reg_3500_pp0_iter1_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter2_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter3_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter4_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter5_reg;
reg   [15:0] mult_386_V_reg_3539;
reg   [15:0] mult_386_V_reg_3539_pp0_iter1_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter2_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter3_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter4_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter5_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter6_reg;
reg   [15:0] mult_449_V_reg_3582;
reg   [15:0] mult_449_V_reg_3582_pp0_iter1_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter2_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter3_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter4_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter5_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter6_reg;
reg   [15:0] mult_512_V_reg_3629;
reg   [15:0] mult_512_V_reg_3629_pp0_iter1_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter2_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter3_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter4_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter5_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter6_reg;
reg   [15:0] mult_576_V_reg_3674;
reg   [15:0] mult_576_V_reg_3674_pp0_iter1_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter2_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter3_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter4_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter5_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter6_reg;
reg   [15:0] mult_640_V_reg_3716;
reg   [15:0] mult_640_V_reg_3716_pp0_iter1_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter2_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter3_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter4_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter5_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter6_reg;
reg   [15:0] mult_704_V_reg_3765;
reg   [15:0] mult_704_V_reg_3765_pp0_iter1_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter2_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter3_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter4_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter5_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter6_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter7_reg;
reg   [15:0] mult_770_V_reg_3814;
reg   [15:0] mult_770_V_reg_3814_pp0_iter1_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter2_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter3_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter4_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter5_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter6_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter7_reg;
reg   [15:0] mult_832_V_reg_3861;
reg   [15:0] mult_832_V_reg_3861_pp0_iter1_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter2_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter3_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter4_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter5_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter6_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter7_reg;
reg   [15:0] mult_896_V_reg_3909;
reg   [15:0] mult_896_V_reg_3909_pp0_iter1_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter2_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter3_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter4_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter5_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter6_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter7_reg;
reg   [15:0] mult_960_V_reg_3958;
reg   [15:0] mult_960_V_reg_3958_pp0_iter1_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter2_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter3_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter4_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter5_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter6_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter7_reg;
wire   [15:0] add_ln703_fu_242_p2;
reg   [15:0] add_ln703_reg_4010;
reg   [15:0] add_ln703_reg_4010_pp0_iter1_reg;
reg   [15:0] add_ln703_reg_4010_pp0_iter2_reg;
wire   [15:0] sub_ln703_fu_248_p2;
reg   [15:0] sub_ln703_reg_4017;
reg   [15:0] sub_ln703_reg_4017_pp0_iter2_reg;
wire   [15:0] sub_ln703_531_fu_252_p2;
reg   [15:0] sub_ln703_531_reg_4023;
reg   [15:0] sub_ln703_531_reg_4023_pp0_iter2_reg;
wire   [15:0] sub_ln703_534_fu_256_p2;
reg   [15:0] sub_ln703_534_reg_4029;
reg   [15:0] sub_ln703_534_reg_4029_pp0_iter2_reg;
reg   [15:0] sub_ln703_534_reg_4029_pp0_iter3_reg;
reg   [15:0] sub_ln703_534_reg_4029_pp0_iter4_reg;
wire   [15:0] add_ln703_539_fu_260_p2;
reg   [15:0] add_ln703_539_reg_4035;
reg   [15:0] add_ln703_539_reg_4035_pp0_iter2_reg;
reg   [15:0] add_ln703_539_reg_4035_pp0_iter3_reg;
wire   [15:0] sub_ln703_533_fu_264_p2;
reg   [15:0] sub_ln703_533_reg_4042;
reg   [15:0] sub_ln703_533_reg_4042_pp0_iter3_reg;
reg   [15:0] sub_ln703_533_reg_4042_pp0_iter4_reg;
wire   [15:0] sub_ln703_538_fu_268_p2;
reg   [15:0] sub_ln703_538_reg_4048;
reg   [15:0] sub_ln703_538_reg_4048_pp0_iter3_reg;
reg   [15:0] sub_ln703_538_reg_4048_pp0_iter4_reg;
reg   [15:0] sub_ln703_538_reg_4048_pp0_iter5_reg;
wire   [15:0] add_ln703_543_fu_272_p2;
reg   [15:0] add_ln703_543_reg_4054;
reg   [15:0] add_ln703_543_reg_4054_pp0_iter3_reg;
reg   [15:0] add_ln703_543_reg_4054_pp0_iter4_reg;
wire   [15:0] sub_ln703_532_fu_276_p2;
reg   [15:0] sub_ln703_532_reg_4061;
reg   [15:0] sub_ln703_532_reg_4061_pp0_iter4_reg;
wire   [15:0] add_ln703_538_fu_280_p2;
reg   [15:0] add_ln703_538_reg_4067;
reg   [15:0] add_ln703_538_reg_4067_pp0_iter4_reg;
wire   [15:0] sub_ln703_535_fu_284_p2;
reg   [15:0] sub_ln703_535_reg_4073;
reg   [15:0] sub_ln703_535_reg_4073_pp0_iter4_reg;
wire   [15:0] add_ln703_540_fu_288_p2;
reg   [15:0] add_ln703_540_reg_4079;
reg   [15:0] add_ln703_540_reg_4079_pp0_iter4_reg;
wire   [15:0] sub_ln703_537_fu_292_p2;
reg   [15:0] sub_ln703_537_reg_4085;
reg   [15:0] sub_ln703_537_reg_4085_pp0_iter4_reg;
reg   [15:0] sub_ln703_537_reg_4085_pp0_iter5_reg;
wire   [15:0] sub_ln703_543_fu_296_p2;
reg   [15:0] sub_ln703_543_reg_4091;
reg   [15:0] sub_ln703_543_reg_4091_pp0_iter4_reg;
wire   [15:0] sub_ln703_545_fu_300_p2;
reg   [15:0] sub_ln703_545_reg_4097;
reg   [15:0] sub_ln703_545_reg_4097_pp0_iter4_reg;
reg   [15:0] sub_ln703_545_reg_4097_pp0_iter5_reg;
wire   [15:0] add_ln703_549_fu_304_p2;
reg   [15:0] add_ln703_549_reg_4103;
reg   [15:0] add_ln703_549_reg_4103_pp0_iter4_reg;
reg   [15:0] add_ln703_549_reg_4103_pp0_iter5_reg;
wire   [15:0] sub_ln703_540_fu_308_p2;
reg   [15:0] sub_ln703_540_reg_4110;
reg   [15:0] sub_ln703_540_reg_4110_pp0_iter5_reg;
wire   [15:0] add_ln703_544_fu_312_p2;
reg   [15:0] add_ln703_544_reg_4116;
reg   [15:0] add_ln703_544_reg_4116_pp0_iter5_reg;
wire   [15:0] sub_ln703_544_fu_316_p2;
reg   [15:0] sub_ln703_544_reg_4122;
reg   [15:0] sub_ln703_544_reg_4122_pp0_iter5_reg;
wire   [15:0] add_ln703_547_fu_320_p2;
reg   [15:0] add_ln703_547_reg_4128;
wire   [15:0] add_ln703_554_fu_324_p2;
reg   [15:0] add_ln703_554_reg_4134;
reg   [15:0] add_ln703_554_reg_4134_pp0_iter5_reg;
wire   [15:0] sub_ln703_558_fu_328_p2;
reg   [15:0] sub_ln703_558_reg_4140;
reg   [15:0] sub_ln703_558_reg_4140_pp0_iter5_reg;
wire   [15:0] add_ln703_559_fu_332_p2;
reg   [15:0] add_ln703_559_reg_4146;
reg   [15:0] add_ln703_559_reg_4146_pp0_iter5_reg;
wire   [15:0] add_ln703_560_fu_336_p2;
reg   [15:0] add_ln703_560_reg_4153;
reg   [15:0] add_ln703_560_reg_4153_pp0_iter5_reg;
wire   [15:0] sub_ln703_536_fu_340_p2;
reg   [15:0] sub_ln703_536_reg_4159;
wire   [15:0] sub_ln703_539_fu_344_p2;
reg   [15:0] sub_ln703_539_reg_4165;
wire   [15:0] add_ln703_541_fu_348_p2;
reg   [15:0] add_ln703_541_reg_4171;
wire   [15:0] add_ln703_542_fu_352_p2;
reg   [15:0] add_ln703_542_reg_4177;
wire   [15:0] add_ln703_545_fu_364_p2;
reg   [15:0] add_ln703_545_reg_4183;
wire   [15:0] add_ln703_548_fu_368_p2;
reg   [15:0] add_ln703_548_reg_4188;
wire   [15:0] sub_ln703_549_fu_372_p2;
reg   [15:0] sub_ln703_549_reg_4194;
wire   [15:0] sub_ln703_550_fu_376_p2;
reg   [15:0] sub_ln703_550_reg_4200;
wire   [15:0] sub_ln703_551_fu_380_p2;
reg   [15:0] sub_ln703_551_reg_4205;
wire   [15:0] add_ln703_550_fu_384_p2;
reg   [15:0] add_ln703_550_reg_4211;
wire   [15:0] sub_ln703_552_fu_388_p2;
reg   [15:0] sub_ln703_552_reg_4217;
wire   [15:0] add_ln703_551_fu_393_p2;
reg   [15:0] add_ln703_551_reg_4222;
wire   [15:0] sub_ln703_554_fu_398_p2;
reg   [15:0] sub_ln703_554_reg_4228;
wire   [15:0] sub_ln703_557_fu_402_p2;
reg   [15:0] sub_ln703_557_reg_4234;
wire   [15:0] add_ln703_564_fu_406_p2;
reg   [15:0] add_ln703_564_reg_4240;
wire   [15:0] sub_ln703_570_fu_410_p2;
reg   [15:0] sub_ln703_570_reg_4246;
wire   [15:0] sub_ln703_576_fu_414_p2;
reg   [15:0] sub_ln703_576_reg_4252;
reg   [15:0] sub_ln703_576_reg_4252_pp0_iter6_reg;
wire   [15:0] add_ln703_566_fu_418_p2;
reg   [15:0] add_ln703_566_reg_4258;
reg   [15:0] add_ln703_566_reg_4258_pp0_iter6_reg;
wire   [15:0] sub_ln703_584_fu_422_p2;
reg   [15:0] sub_ln703_584_reg_4264;
reg   [15:0] sub_ln703_584_reg_4264_pp0_iter6_reg;
wire   [15:0] add_ln703_568_fu_426_p2;
reg   [15:0] add_ln703_568_reg_4270;
wire   [15:0] sub_ln703_591_fu_430_p2;
reg   [15:0] sub_ln703_591_reg_4277;
wire   [15:0] add_ln703_597_fu_434_p2;
reg   [15:0] add_ln703_597_reg_4282;
reg   [15:0] add_ln703_597_reg_4282_pp0_iter6_reg;
wire   [15:0] add_ln703_557_fu_488_p2;
reg   [15:0] add_ln703_557_reg_4293;
wire   [15:0] add_ln703_558_fu_498_p2;
reg   [15:0] add_ln703_558_reg_4298;
wire   [15:0] sub_ln703_567_fu_540_p2;
reg   [15:0] sub_ln703_567_reg_4303;
wire   [15:0] sub_ln703_572_fu_563_p2;
reg   [15:0] sub_ln703_572_reg_4309;
wire   [15:0] sub_ln703_574_fu_572_p2;
reg   [15:0] sub_ln703_574_reg_4314;
wire   [15:0] sub_ln703_578_fu_585_p2;
reg   [15:0] sub_ln703_578_reg_4319;
wire   [15:0] sub_ln703_579_fu_590_p2;
reg   [15:0] sub_ln703_579_reg_4324;
wire   [15:0] sub_ln703_582_fu_599_p2;
reg   [15:0] sub_ln703_582_reg_4329;
wire   [15:0] sub_ln703_585_fu_609_p2;
reg   [15:0] sub_ln703_585_reg_4334;
wire   [15:0] sub_ln703_586_fu_614_p2;
reg   [15:0] sub_ln703_586_reg_4340;
wire   [15:0] sub_ln703_587_fu_619_p2;
reg   [15:0] sub_ln703_587_reg_4345;
wire   [15:0] sub_ln703_588_fu_624_p2;
reg   [15:0] sub_ln703_588_reg_4350;
wire   [15:0] sub_ln703_589_fu_638_p2;
reg   [15:0] sub_ln703_589_reg_4355;
wire   [15:0] sub_ln703_590_fu_643_p2;
reg   [15:0] sub_ln703_590_reg_4361;
wire   [15:0] sub_ln703_592_fu_653_p2;
reg   [15:0] sub_ln703_592_reg_4366;
wire   [15:0] add_ln703_571_fu_657_p2;
reg   [15:0] add_ln703_571_reg_4372;
wire   [15:0] sub_ln703_594_fu_666_p2;
reg   [15:0] sub_ln703_594_reg_4377;
wire   [15:0] add_ln703_572_fu_670_p2;
reg   [15:0] add_ln703_572_reg_4382;
wire   [15:0] add_ln703_573_fu_675_p2;
reg   [15:0] add_ln703_573_reg_4387;
wire   [15:0] add_ln703_574_fu_679_p2;
reg   [15:0] add_ln703_574_reg_4393;
wire   [15:0] sub_ln703_596_fu_683_p2;
reg   [15:0] sub_ln703_596_reg_4398;
wire   [15:0] sub_ln703_599_fu_693_p2;
reg   [15:0] sub_ln703_599_reg_4403;
wire   [15:0] add_ln703_576_fu_702_p2;
reg   [15:0] add_ln703_576_reg_4408;
wire   [15:0] add_ln703_577_fu_707_p2;
reg   [15:0] add_ln703_577_reg_4413;
wire   [15:0] add_ln703_579_fu_716_p2;
reg   [15:0] add_ln703_579_reg_4418;
wire   [15:0] sub_ln703_605_fu_720_p2;
reg   [15:0] sub_ln703_605_reg_4423;
wire   [15:0] sub_ln703_608_fu_725_p2;
reg   [15:0] sub_ln703_608_reg_4428;
wire   [15:0] add_ln703_580_fu_730_p2;
reg   [15:0] add_ln703_580_reg_4433;
wire   [15:0] sub_ln703_610_fu_734_p2;
reg   [15:0] sub_ln703_610_reg_4439;
wire   [15:0] sub_ln703_611_fu_739_p2;
reg   [15:0] sub_ln703_611_reg_4444;
wire   [15:0] add_ln703_583_fu_754_p2;
reg   [15:0] add_ln703_583_reg_4450;
wire   [15:0] sub_ln703_613_fu_758_p2;
reg   [15:0] sub_ln703_613_reg_4455;
wire   [15:0] sub_ln703_617_fu_763_p2;
reg   [15:0] sub_ln703_617_reg_4460;
wire   [15:0] sub_ln703_620_fu_772_p2;
reg   [15:0] sub_ln703_620_reg_4466;
wire   [15:0] add_ln703_587_fu_786_p2;
reg   [15:0] add_ln703_587_reg_4471;
wire   [15:0] add_ln703_588_fu_792_p2;
reg   [15:0] add_ln703_588_reg_4476;
wire   [15:0] add_ln703_590_fu_801_p2;
reg   [15:0] add_ln703_590_reg_4481;
wire   [15:0] sub_ln703_627_fu_807_p2;
reg   [15:0] sub_ln703_627_reg_4486;
wire   [15:0] sub_ln703_632_fu_818_p2;
reg   [15:0] sub_ln703_632_reg_4491;
wire   [15:0] sub_ln703_641_fu_838_p2;
reg   [15:0] sub_ln703_641_reg_4496;
wire   [15:0] sub_ln703_645_fu_843_p2;
reg   [15:0] sub_ln703_645_reg_4501;
wire   [15:0] sub_ln703_660_fu_872_p2;
reg   [15:0] sub_ln703_660_reg_4506;
wire   [15:0] sub_ln703_661_fu_877_p2;
reg   [15:0] sub_ln703_661_reg_4511;
wire   [15:0] sub_ln703_662_fu_882_p2;
reg   [15:0] sub_ln703_662_reg_4516;
wire   [15:0] add_ln703_611_fu_887_p2;
reg   [15:0] add_ln703_611_reg_4521;
wire   [15:0] add_ln703_620_fu_891_p2;
reg   [15:0] add_ln703_620_reg_4537;
wire   [15:0] sub_ln703_671_fu_896_p2;
reg   [15:0] sub_ln703_671_reg_4543;
wire   [15:0] sub_ln703_676_fu_901_p2;
reg   [15:0] sub_ln703_676_reg_4548;
wire   [15:0] add_ln703_637_fu_906_p2;
reg   [15:0] add_ln703_637_reg_4553;
wire   [15:0] add_ln703_655_fu_910_p2;
reg   [15:0] add_ln703_655_reg_4558;
wire   [15:0] add_ln703_659_fu_914_p2;
reg   [15:0] add_ln703_659_reg_4568;
wire   [15:0] add_ln703_692_fu_920_p2;
reg   [15:0] add_ln703_692_reg_4573;
reg   [15:0] add_ln703_692_reg_4573_pp0_iter7_reg;
wire   [15:0] add_ln703_631_fu_1397_p2;
reg   [15:0] add_ln703_631_reg_4588;
wire   [15:0] add_ln703_634_fu_1416_p2;
reg   [15:0] add_ln703_634_reg_4593;
wire   [15:0] sub_ln703_692_fu_1433_p2;
reg   [15:0] sub_ln703_692_reg_4598;
wire   [15:0] sub_ln703_693_fu_1438_p2;
reg   [15:0] sub_ln703_693_reg_4603;
wire   [15:0] add_ln703_639_fu_1459_p2;
reg   [15:0] add_ln703_639_reg_4608;
wire   [15:0] sub_ln703_695_fu_1464_p2;
reg   [15:0] sub_ln703_695_reg_4613;
wire   [15:0] sub_ln703_699_fu_1495_p2;
reg   [15:0] sub_ln703_699_reg_4618;
wire   [15:0] sub_ln703_700_fu_1500_p2;
reg   [15:0] sub_ln703_700_reg_4623;
wire   [15:0] add_ln703_642_fu_1505_p2;
reg   [15:0] add_ln703_642_reg_4628;
wire   [15:0] sub_ln703_701_fu_1509_p2;
reg   [15:0] sub_ln703_701_reg_4633;
wire   [15:0] sub_ln703_702_fu_1514_p2;
reg   [15:0] sub_ln703_702_reg_4638;
wire   [15:0] sub_ln703_704_fu_1524_p2;
reg   [15:0] sub_ln703_704_reg_4643;
wire   [15:0] add_ln703_645_fu_1538_p2;
reg   [15:0] add_ln703_645_reg_4648;
wire   [15:0] sub_ln703_706_fu_1548_p2;
reg   [15:0] sub_ln703_706_reg_4653;
wire   [15:0] add_ln703_646_fu_1553_p2;
reg   [15:0] add_ln703_646_reg_4658;
wire   [15:0] sub_ln703_707_fu_1559_p2;
reg   [15:0] sub_ln703_707_reg_4663;
wire   [15:0] sub_ln703_708_fu_1564_p2;
reg   [15:0] sub_ln703_708_reg_4668;
wire   [15:0] sub_ln703_709_fu_1569_p2;
reg   [15:0] sub_ln703_709_reg_4673;
wire   [15:0] sub_ln703_710_fu_1606_p2;
reg   [15:0] sub_ln703_710_reg_4678;
wire   [15:0] sub_ln703_711_fu_1611_p2;
reg   [15:0] sub_ln703_711_reg_4683;
wire   [15:0] sub_ln703_712_fu_1616_p2;
reg   [15:0] sub_ln703_712_reg_4688;
wire   [15:0] sub_ln703_714_fu_1626_p2;
reg   [15:0] sub_ln703_714_reg_4693;
wire   [15:0] sub_ln703_715_fu_1631_p2;
reg   [15:0] sub_ln703_715_reg_4698;
wire   [15:0] sub_ln703_716_fu_1636_p2;
reg   [15:0] sub_ln703_716_reg_4703;
wire   [15:0] sub_ln703_718_fu_1646_p2;
reg   [15:0] sub_ln703_718_reg_4708;
wire   [15:0] sub_ln703_720_fu_1676_p2;
reg   [15:0] sub_ln703_720_reg_4713;
wire   [15:0] sub_ln703_722_fu_1681_p2;
reg   [15:0] sub_ln703_722_reg_4718;
wire   [15:0] sub_ln703_724_fu_1686_p2;
reg   [15:0] sub_ln703_724_reg_4723;
wire   [15:0] sub_ln703_725_fu_1691_p2;
reg   [15:0] sub_ln703_725_reg_4728;
wire   [15:0] add_ln703_658_fu_1696_p2;
reg   [15:0] add_ln703_658_reg_4733;
wire   [15:0] sub_ln703_727_fu_1701_p2;
reg   [15:0] sub_ln703_727_reg_4738;
wire   [15:0] add_ln703_661_fu_1710_p2;
reg   [15:0] add_ln703_661_reg_4744;
wire   [15:0] sub_ln703_729_fu_1715_p2;
reg   [15:0] sub_ln703_729_reg_4749;
wire   [15:0] sub_ln703_730_fu_1720_p2;
reg   [15:0] sub_ln703_730_reg_4754;
wire   [15:0] sub_ln703_731_fu_1725_p2;
reg   [15:0] sub_ln703_731_reg_4759;
wire   [15:0] add_ln703_663_fu_1735_p2;
reg   [15:0] add_ln703_663_reg_4764;
wire   [15:0] sub_ln703_732_fu_1741_p2;
reg   [15:0] sub_ln703_732_reg_4769;
wire   [15:0] sub_ln703_738_fu_1757_p2;
reg   [15:0] sub_ln703_738_reg_4774;
wire   [15:0] sub_ln703_742_fu_1762_p2;
reg   [15:0] sub_ln703_742_reg_4779;
wire   [15:0] add_ln703_667_fu_1767_p2;
reg   [15:0] add_ln703_667_reg_4784;
wire   [15:0] sub_ln703_743_fu_1772_p2;
reg   [15:0] sub_ln703_743_reg_4789;
wire   [15:0] sub_ln703_744_fu_1777_p2;
reg   [15:0] sub_ln703_744_reg_4794;
wire   [15:0] sub_ln703_745_fu_1782_p2;
reg   [15:0] sub_ln703_745_reg_4799;
wire   [15:0] add_ln703_669_fu_1787_p2;
reg   [15:0] add_ln703_669_reg_4804;
wire   [15:0] sub_ln703_748_fu_1792_p2;
reg   [15:0] sub_ln703_748_reg_4809;
wire   [15:0] sub_ln703_751_fu_1797_p2;
reg   [15:0] sub_ln703_751_reg_4814;
wire   [15:0] add_ln703_670_fu_1802_p2;
reg   [15:0] add_ln703_670_reg_4819;
wire   [15:0] sub_ln703_752_fu_1807_p2;
reg   [15:0] sub_ln703_752_reg_4824;
wire   [15:0] add_ln703_672_fu_1812_p2;
reg   [15:0] add_ln703_672_reg_4829;
wire   [15:0] sub_ln703_753_fu_1817_p2;
reg   [15:0] sub_ln703_753_reg_4834;
wire   [15:0] add_ln703_674_fu_1822_p2;
reg   [15:0] add_ln703_674_reg_4839;
wire   [15:0] add_ln703_679_fu_1826_p2;
reg   [15:0] add_ln703_679_reg_4847;
wire   [15:0] sub_ln703_765_fu_1832_p2;
reg   [15:0] sub_ln703_765_reg_4852;
wire   [15:0] add_ln703_687_fu_1847_p2;
reg   [15:0] add_ln703_687_reg_4857;
wire   [15:0] add_ln703_688_fu_1853_p2;
reg   [15:0] add_ln703_688_reg_4862;
wire   [15:0] add_ln703_707_fu_1877_p2;
reg   [15:0] add_ln703_707_reg_4867;
wire   [15:0] add_ln703_711_fu_1887_p2;
reg   [15:0] add_ln703_711_reg_4872;
wire   [15:0] add_ln703_716_fu_1902_p2;
reg   [15:0] add_ln703_716_reg_4877;
wire   [15:0] add_ln703_722_fu_1913_p2;
reg   [15:0] add_ln703_722_reg_4882;
wire   [15:0] add_ln703_724_fu_1923_p2;
reg   [15:0] add_ln703_724_reg_4887;
wire   [15:0] add_ln703_727_fu_1934_p2;
reg   [15:0] add_ln703_727_reg_4892;
wire   [15:0] add_ln703_729_fu_1945_p2;
reg   [15:0] add_ln703_729_reg_4897;
wire   [15:0] add_ln703_732_fu_1956_p2;
reg   [15:0] add_ln703_732_reg_4902;
wire   [15:0] add_ln703_737_fu_1962_p2;
reg   [15:0] add_ln703_737_reg_4907;
wire   [15:0] add_ln703_739_fu_1966_p2;
reg   [15:0] add_ln703_739_reg_4915;
wire   [15:0] add_ln703_751_fu_1971_p2;
reg   [15:0] add_ln703_751_reg_4920;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_541_fu_356_p2;
wire   [15:0] sub_ln703_542_fu_360_p2;
wire   [15:0] add_ln703_546_fu_438_p2;
wire   [15:0] sub_ln703_546_fu_442_p2;
wire   [15:0] sub_ln703_547_fu_446_p2;
wire   [15:0] sub_ln703_548_fu_450_p2;
wire   [15:0] add_ln703_552_fu_454_p2;
wire   [15:0] add_ln703_553_fu_458_p2;
wire   [15:0] sub_ln703_553_fu_462_p2;
wire   [15:0] add_ln703_555_fu_466_p2;
wire   [15:0] sub_ln703_555_fu_470_p2;
wire   [15:0] sub_ln703_556_fu_474_p2;
wire   [15:0] add_ln703_556_fu_478_p2;
wire   [15:0] sub_ln703_559_fu_483_p2;
wire   [15:0] sub_ln703_560_fu_493_p2;
wire   [15:0] sub_ln703_561_fu_502_p2;
wire   [15:0] sub_ln703_562_fu_506_p2;
wire   [15:0] add_ln703_561_fu_510_p2;
wire   [15:0] add_ln703_562_fu_522_p2;
wire   [15:0] add_ln703_567_fu_629_p2;
wire   [15:0] add_ln703_563_fu_526_p2;
wire   [15:0] sub_ln703_565_fu_530_p2;
wire   [15:0] sub_ln703_566_fu_535_p2;
wire   [15:0] sub_ln703_568_fu_545_p2;
wire   [15:0] sub_ln703_569_fu_549_p2;
wire   [15:0] add_ln703_565_fu_554_p2;
wire   [15:0] sub_ln703_571_fu_558_p2;
wire   [15:0] sub_ln703_573_fu_567_p2;
wire   [15:0] sub_ln703_575_fu_577_p2;
wire   [15:0] sub_ln703_577_fu_581_p2;
wire   [15:0] sub_ln703_580_fu_594_p2;
wire   [15:0] sub_ln703_583_fu_604_p2;
wire   [15:0] sub_ln703_564_fu_518_p2;
wire   [15:0] add_ln703_581_fu_744_p2;
wire   [15:0] add_ln703_569_fu_633_p2;
wire   [15:0] add_ln703_570_fu_648_p2;
wire   [15:0] sub_ln703_593_fu_661_p2;
wire   [15:0] add_ln703_585_fu_777_p2;
wire   [15:0] add_ln703_586_fu_781_p2;
wire   [15:0] sub_ln703_597_fu_688_p2;
wire   [15:0] add_ln703_589_fu_797_p2;
wire   [15:0] add_ln703_575_fu_698_p2;
wire   [15:0] sub_ln703_602_fu_712_p2;
wire   [15:0] add_ln703_595_fu_828_p2;
wire   [15:0] add_ln703_582_fu_748_p2;
wire   [15:0] sub_ln703_618_fu_768_p2;
wire   [15:0] add_ln703_600_fu_848_p2;
wire   [15:0] add_ln703_601_fu_852_p2;
wire   [15:0] add_ln703_605_fu_862_p2;
wire   [15:0] add_ln703_593_fu_812_p2;
wire   [15:0] add_ln703_594_fu_823_p2;
wire   [15:0] add_ln703_596_fu_832_p2;
wire   [15:0] add_ln703_602_fu_856_p2;
wire   [15:0] add_ln703_606_fu_866_p2;
wire   [15:0] sub_ln703_563_fu_514_p2;
wire   [15:0] sub_ln703_581_fu_924_p2;
wire   [15:0] sub_ln703_595_fu_928_p2;
wire   [15:0] sub_ln703_600_fu_936_p2;
wire   [15:0] add_ln703_578_fu_944_p2;
wire   [15:0] sub_ln703_607_fu_961_p2;
wire   [15:0] sub_ln703_609_fu_965_p2;
wire   [15:0] sub_ln703_612_fu_969_p2;
wire   [15:0] add_ln703_584_fu_985_p2;
wire   [15:0] sub_ln703_621_fu_993_p2;
wire   [15:0] sub_ln703_623_fu_1002_p2;
wire   [15:0] sub_ln703_624_fu_1006_p2;
wire   [15:0] sub_ln703_625_fu_1010_p2;
wire   [15:0] sub_ln703_598_fu_932_p2;
wire   [15:0] add_ln703_591_fu_1027_p2;
wire   [15:0] add_ln703_592_fu_1031_p2;
wire   [15:0] sub_ln703_630_fu_1035_p2;
wire   [15:0] sub_ln703_631_fu_1039_p2;
wire   [15:0] add_ln703_598_fu_1052_p2;
wire   [15:0] sub_ln703_604_fu_952_p2;
wire   [15:0] sub_ln703_635_fu_1056_p2;
wire   [15:0] sub_ln703_637_fu_1065_p2;
wire   [15:0] sub_ln703_638_fu_1069_p2;
wire   [15:0] add_ln703_599_fu_1073_p2;
wire   [15:0] sub_ln703_639_fu_1078_p2;
wire   [15:0] sub_ln703_643_fu_1091_p2;
wire   [15:0] sub_ln703_644_fu_1095_p2;
wire   [15:0] sub_ln703_615_fu_977_p2;
wire   [15:0] sub_ln703_616_fu_981_p2;
wire   [15:0] sub_ln703_646_fu_1099_p2;
wire   [15:0] sub_ln703_636_fu_1060_p2;
wire   [15:0] sub_ln703_647_fu_1104_p2;
wire   [15:0] sub_ln703_648_fu_1108_p2;
wire   [15:0] sub_ln703_649_fu_1113_p2;
wire   [15:0] sub_ln703_651_fu_1122_p2;
wire   [15:0] sub_ln703_652_fu_1127_p2;
wire   [15:0] add_ln703_603_fu_1132_p2;
wire   [15:0] sub_ln703_653_fu_1136_p2;
wire   [15:0] add_ln703_604_fu_1140_p2;
wire   [15:0] sub_ln703_655_fu_1149_p2;
wire   [15:0] sub_ln703_629_fu_1022_p2;
wire   [15:0] sub_ln703_656_fu_1153_p2;
wire   [15:0] add_ln703_626_fu_1321_p2;
wire   [15:0] sub_ln703_657_fu_1158_p2;
wire   [15:0] add_ln703_607_fu_1163_p2;
wire   [15:0] sub_ln703_658_fu_1167_p2;
wire   [15:0] sub_ln703_659_fu_1171_p2;
wire   [15:0] sub_ln703_601_fu_940_p2;
wire   [15:0] add_ln703_628_fu_1350_p2;
wire   [15:0] add_ln703_608_fu_1176_p2;
wire   [15:0] add_ln703_609_fu_1181_p2;
wire   [15:0] add_ln703_610_fu_1185_p2;
wire   [15:0] sub_ln703_634_fu_1048_p2;
wire   [15:0] sub_ln703_663_fu_1189_p2;
wire   [15:0] add_ln703_612_fu_1194_p2;
wire   [15:0] sub_ln703_664_fu_1199_p2;
wire   [15:0] sub_ln703_606_fu_956_p2;
wire   [15:0] add_ln703_632_fu_1407_p2;
wire   [15:0] add_ln703_633_fu_1412_p2;
wire   [15:0] sub_ln703_665_fu_1204_p2;
wire   [15:0] add_ln703_613_fu_1209_p2;
wire   [15:0] sub_ln703_666_fu_1214_p2;
wire   [15:0] add_ln703_614_fu_1219_p2;
wire   [15:0] sub_ln703_640_fu_1082_p2;
wire   [15:0] add_ln703_638_fu_1454_p2;
wire   [15:0] sub_ln703_667_fu_1224_p2;
wire   [15:0] sub_ln703_642_fu_1086_p2;
wire   [15:0] add_ln703_615_fu_1228_p2;
wire   [15:0] sub_ln703_668_fu_1233_p2;
wire   [15:0] add_ln703_616_fu_1238_p2;
wire   [15:0] add_ln703_617_fu_1243_p2;
wire   [15:0] add_ln703_618_fu_1248_p2;
wire   [15:0] add_ln703_619_fu_1252_p2;
wire   [15:0] add_ln703_621_fu_1256_p2;
wire   [15:0] sub_ln703_669_fu_1261_p2;
wire   [15:0] sub_ln703_670_fu_1266_p2;
wire   [15:0] add_ln703_622_fu_1271_p2;
wire   [15:0] add_ln703_643_fu_1529_p2;
wire   [15:0] add_ln703_644_fu_1533_p2;
wire   [15:0] add_ln703_623_fu_1276_p2;
wire   [15:0] sub_ln703_650_fu_1118_p2;
wire   [15:0] sub_ln703_672_fu_1281_p2;
wire   [15:0] add_ln703_624_fu_1286_p2;
wire   [15:0] sub_ln703_674_fu_1296_p2;
wire   [15:0] sub_ln703_626_fu_1014_p2;
wire   [15:0] add_ln703_648_fu_1579_p2;
wire   [15:0] sub_ln703_677_fu_1306_p2;
wire   [15:0] sub_ln703_628_fu_1018_p2;
wire   [15:0] add_ln703_651_fu_1595_p2;
wire   [15:0] add_ln703_625_fu_1311_p2;
wire   [15:0] sub_ln703_678_fu_1316_p2;
wire   [15:0] add_ln703_627_fu_1325_p2;
wire   [15:0] sub_ln703_681_fu_1340_p2;
wire   [15:0] sub_ln703_682_fu_1345_p2;
wire   [15:0] add_ln703_629_fu_1355_p2;
wire   [15:0] sub_ln703_683_fu_1360_p2;
wire   [15:0] sub_ln703_684_fu_1365_p2;
wire   [15:0] sub_ln703_686_fu_1374_p2;
wire   [15:0] sub_ln703_687_fu_1378_p2;
wire   [15:0] add_ln703_630_fu_1387_p2;
wire   [15:0] sub_ln703_603_fu_948_p2;
wire   [15:0] add_ln703_654_fu_1661_p2;
wire   [15:0] add_ln703_656_fu_1666_p2;
wire   [15:0] sub_ln703_689_fu_1392_p2;
wire   [15:0] sub_ln703_690_fu_1402_p2;
wire   [15:0] add_ln703_635_fu_1422_p2;
wire   [15:0] sub_ln703_691_fu_1428_p2;
wire   [15:0] sub_ln703_694_fu_1443_p2;
wire   [15:0] add_ln703_636_fu_1448_p2;
wire   [15:0] add_ln703_660_fu_1706_p2;
wire   [15:0] add_ln703_640_fu_1469_p2;
wire   [15:0] sub_ln703_696_fu_1475_p2;
wire   [15:0] add_ln703_641_fu_1480_p2;
wire   [15:0] sub_ln703_614_fu_973_p2;
wire   [15:0] add_ln703_662_fu_1730_p2;
wire   [15:0] sub_ln703_697_fu_1485_p2;
wire   [15:0] sub_ln703_619_fu_989_p2;
wire   [15:0] add_ln703_665_fu_1746_p2;
wire   [15:0] sub_ln703_705_fu_1544_p2;
wire   [15:0] add_ln703_647_fu_1574_p2;
wire   [15:0] sub_ln703_675_fu_1301_p2;
wire   [15:0] add_ln703_649_fu_1584_p2;
wire   [15:0] add_ln703_650_fu_1590_p2;
wire   [15:0] add_ln703_652_fu_1600_p2;
wire   [15:0] sub_ln703_680_fu_1335_p2;
wire   [15:0] sub_ln703_713_fu_1621_p2;
wire   [15:0] sub_ln703_717_fu_1641_p2;
wire   [15:0] sub_ln703_685_fu_1370_p2;
wire   [15:0] add_ln703_653_fu_1651_p2;
wire   [15:0] sub_ln703_719_fu_1656_p2;
wire   [15:0] add_ln703_657_fu_1670_p2;
wire   [15:0] sub_ln703_698_fu_1490_p2;
wire   [15:0] add_ln703_666_fu_1751_p2;
wire   [15:0] sub_ln703_654_fu_1145_p2;
wire   [15:0] add_ln703_685_fu_1837_p2;
wire   [15:0] add_ln703_686_fu_1842_p2;
wire   [15:0] sub_ln703_679_fu_1330_p2;
wire   [15:0] add_ln703_703_fu_1858_p2;
wire   [15:0] add_ln703_705_fu_1867_p2;
wire   [15:0] add_ln703_704_fu_1862_p2;
wire   [15:0] add_ln703_706_fu_1871_p2;
wire   [15:0] add_ln703_710_fu_1883_p2;
wire   [15:0] sub_ln703_622_fu_997_p2;
wire   [15:0] add_ln703_714_fu_1893_p2;
wire   [15:0] add_ln703_715_fu_1898_p2;
wire   [15:0] sub_ln703_673_fu_1291_p2;
wire   [15:0] add_ln703_721_fu_1908_p2;
wire   [15:0] add_ln703_723_fu_1919_p2;
wire   [15:0] add_ln703_726_fu_1929_p2;
wire   [15:0] sub_ln703_633_fu_1043_p2;
wire   [15:0] add_ln703_728_fu_1940_p2;
wire   [15:0] sub_ln703_688_fu_1382_p2;
wire   [15:0] add_ln703_731_fu_1951_p2;
wire   [15:0] sub_ln703_703_fu_1519_p2;
wire   [15:0] sub_ln703_723_fu_1979_p2;
wire   [15:0] sub_ln703_726_fu_1983_p2;
wire   [15:0] add_ln703_664_fu_1991_p2;
wire   [15:0] sub_ln703_736_fu_2007_p2;
wire   [15:0] sub_ln703_739_fu_2015_p2;
wire   [15:0] sub_ln703_740_fu_2019_p2;
wire   [15:0] sub_ln703_741_fu_2023_p2;
wire   [15:0] sub_ln703_746_fu_2027_p2;
wire   [15:0] sub_ln703_747_fu_2031_p2;
wire   [15:0] add_ln703_668_fu_2035_p2;
wire   [15:0] sub_ln703_749_fu_2039_p2;
wire   [15:0] sub_ln703_750_fu_2043_p2;
wire   [15:0] add_ln703_671_fu_2047_p2;
wire   [15:0] sub_ln703_754_fu_2051_p2;
wire   [15:0] sub_ln703_721_fu_1975_p2;
wire   [15:0] sub_ln703_755_fu_2055_p2;
wire   [15:0] sub_ln703_757_fu_2064_p2;
wire   [15:0] add_ln703_673_fu_2068_p2;
wire   [15:0] add_ln703_675_fu_2072_p2;
wire   [15:0] sub_ln703_758_fu_2076_p2;
wire   [15:0] sub_ln703_759_fu_2081_p2;
wire   [15:0] sub_ln703_728_fu_1987_p2;
wire   [15:0] sub_ln703_761_fu_2089_p2;
wire   [15:0] add_ln703_676_fu_2093_p2;
wire   [15:0] sub_ln703_762_fu_2097_p2;
wire   [15:0] add_ln703_677_fu_2101_p2;
wire   [15:0] sub_ln703_763_fu_2105_p2;
wire   [15:0] add_ln703_678_fu_2109_p2;
wire   [15:0] sub_ln703_733_fu_1995_p2;
wire   [15:0] sub_ln703_734_fu_1999_p2;
wire   [15:0] sub_ln703_735_fu_2003_p2;
wire   [15:0] add_ln703_680_fu_2118_p2;
wire   [15:0] add_ln703_708_fu_2323_p2;
wire   [15:0] sub_ln703_737_fu_2011_p2;
wire   [15:0] sub_ln703_766_fu_2123_p2;
wire   [15:0] add_ln703_717_fu_2342_p2;
wire   [15:0] add_ln703_681_fu_2132_p2;
wire   [15:0] add_ln703_682_fu_2136_p2;
wire   [15:0] add_ln703_719_fu_2361_p2;
wire   [15:0] add_ln703_683_fu_2146_p2;
wire   [15:0] sub_ln703_769_fu_2150_p2;
wire   [15:0] add_ln703_684_fu_2154_p2;
wire   [15:0] sub_ln703_770_fu_2158_p2;
wire   [15:0] sub_ln703_771_fu_2162_p2;
wire   [15:0] add_ln703_689_fu_2181_p2;
wire   [15:0] sub_ln703_775_fu_2185_p2;
wire   [15:0] add_ln703_690_fu_2189_p2;
wire   [15:0] add_ln703_691_fu_2193_p2;
wire   [15:0] sub_ln703_778_fu_2207_p2;
wire   [15:0] sub_ln703_779_fu_2211_p2;
wire   [15:0] sub_ln703_780_fu_2215_p2;
wire   [15:0] sub_ln703_781_fu_2220_p2;
wire   [15:0] sub_ln703_782_fu_2224_p2;
wire   [15:0] add_ln703_693_fu_2229_p2;
wire   [15:0] add_ln703_694_fu_2234_p2;
wire   [15:0] add_ln703_695_fu_2239_p2;
wire   [15:0] sub_ln703_783_fu_2244_p2;
wire   [15:0] sub_ln703_784_fu_2249_p2;
wire   [15:0] sub_ln703_786_fu_2259_p2;
wire   [15:0] add_ln703_696_fu_2264_p2;
wire   [15:0] add_ln703_697_fu_2269_p2;
wire   [15:0] sub_ln703_787_fu_2274_p2;
wire   [15:0] add_ln703_698_fu_2279_p2;
wire   [15:0] sub_ln703_788_fu_2284_p2;
wire   [15:0] add_ln703_699_fu_2289_p2;
wire   [15:0] sub_ln703_789_fu_2294_p2;
wire   [15:0] add_ln703_700_fu_2303_p2;
wire   [15:0] add_ln703_701_fu_2308_p2;
wire   [15:0] add_ln703_702_fu_2313_p2;
wire   [15:0] add_ln703_740_fu_2532_p2;
wire   [15:0] add_ln703_709_fu_2327_p2;
wire   [15:0] add_ln703_712_fu_2332_p2;
wire   [15:0] add_ln703_713_fu_2337_p2;
wire   [15:0] add_ln703_718_fu_2346_p2;
wire   [15:0] sub_ln703_792_fu_2351_p2;
wire   [15:0] add_ln703_720_fu_2365_p2;
wire   [15:0] sub_ln703_768_fu_2141_p2;
wire   [15:0] sub_ln703_794_fu_2370_p2;
wire   [15:0] sub_ln703_795_fu_2375_p2;
wire   [15:0] sub_ln703_796_fu_2380_p2;
wire   [15:0] add_ln703_725_fu_2389_p2;
wire   [15:0] sub_ln703_798_fu_2394_p2;
wire   [15:0] sub_ln703_799_fu_2399_p2;
wire   [15:0] sub_ln703_800_fu_2404_p2;
wire   [15:0] sub_ln703_801_fu_2409_p2;
wire   [15:0] sub_ln703_802_fu_2414_p2;
wire   [15:0] sub_ln703_776_fu_2197_p2;
wire   [15:0] sub_ln703_803_fu_2419_p2;
wire   [15:0] add_ln703_730_fu_2424_p2;
wire   [15:0] add_ln703_733_fu_2434_p2;
wire   [15:0] add_ln703_750_fu_2669_p2;
wire   [15:0] sub_ln703_805_fu_2439_p2;
wire   [15:0] sub_ln703_806_fu_2444_p2;
wire   [15:0] sub_ln703_807_fu_2449_p2;
wire   [15:0] sub_ln703_756_fu_2059_p2;
wire   [15:0] add_ln703_754_fu_2693_p2;
wire   [15:0] sub_ln703_808_fu_2454_p2;
wire   [15:0] sub_ln703_809_fu_2459_p2;
wire   [15:0] sub_ln703_810_fu_2464_p2;
wire   [15:0] sub_ln703_785_fu_2254_p2;
wire   [15:0] add_ln703_734_fu_2469_p2;
wire   [15:0] sub_ln703_760_fu_2085_p2;
wire   [15:0] add_ln703_758_fu_2728_p2;
wire   [15:0] sub_ln703_811_fu_2474_p2;
wire   [15:0] sub_ln703_812_fu_2479_p2;
wire   [15:0] add_ln703_735_fu_2484_p2;
wire   [15:0] sub_ln703_813_fu_2489_p2;
wire   [15:0] sub_ln703_814_fu_2494_p2;
wire   [15:0] add_ln703_761_fu_2763_p2;
wire   [15:0] add_ln703_762_fu_2767_p2;
wire   [15:0] sub_ln703_815_fu_2499_p2;
wire   [15:0] add_ln703_736_fu_2504_p2;
wire   [15:0] sub_ln703_790_fu_2299_p2;
wire   [15:0] sub_ln703_764_fu_2113_p2;
wire   [15:0] add_ln703_765_fu_2792_p2;
wire   [15:0] sub_ln703_816_fu_2509_p2;
wire   [15:0] sub_ln703_817_fu_2514_p2;
wire   [15:0] sub_ln703_818_fu_2519_p2;
wire   [15:0] sub_ln703_819_fu_2524_p2;
wire   [15:0] sub_ln703_791_fu_2318_p2;
wire   [15:0] add_ln703_738_fu_2528_p2;
wire   [15:0] add_ln703_741_fu_2536_p2;
wire   [15:0] sub_ln703_820_fu_2541_p2;
wire   [15:0] sub_ln703_821_fu_2546_p2;
wire   [15:0] sub_ln703_822_fu_2550_p2;
wire   [15:0] sub_ln703_823_fu_2555_p2;
wire   [15:0] sub_ln703_824_fu_2560_p2;
wire   [15:0] sub_ln703_825_fu_2564_p2;
wire   [15:0] sub_ln703_767_fu_2127_p2;
wire   [15:0] add_ln703_770_fu_2867_p2;
wire   [15:0] add_ln703_742_fu_2569_p2;
wire   [15:0] sub_ln703_793_fu_2356_p2;
wire   [15:0] sub_ln703_826_fu_2574_p2;
wire   [15:0] sub_ln703_827_fu_2579_p2;
wire   [15:0] add_ln703_743_fu_2583_p2;
wire   [15:0] sub_ln703_828_fu_2588_p2;
wire   [15:0] sub_ln703_829_fu_2593_p2;
wire   [15:0] sub_ln703_830_fu_2598_p2;
wire   [15:0] sub_ln703_831_fu_2602_p2;
wire   [15:0] sub_ln703_797_fu_2385_p2;
wire   [15:0] sub_ln703_832_fu_2607_p2;
wire   [15:0] add_ln703_744_fu_2612_p2;
wire   [15:0] sub_ln703_772_fu_2166_p2;
wire   [15:0] add_ln703_776_fu_2937_p2;
wire   [15:0] sub_ln703_773_fu_2171_p2;
wire   [15:0] add_ln703_778_fu_2947_p2;
wire   [15:0] sub_ln703_774_fu_2176_p2;
wire   [15:0] add_ln703_780_fu_2957_p2;
wire   [15:0] add_ln703_745_fu_2617_p2;
wire   [15:0] add_ln703_746_fu_2622_p2;
wire   [15:0] add_ln703_747_fu_2627_p2;
wire   [15:0] add_ln703_748_fu_2632_p2;
wire   [15:0] add_ln703_749_fu_2637_p2;
wire   [15:0] sub_ln703_777_fu_2202_p2;
wire   [15:0] add_ln703_782_fu_2992_p2;
wire   [15:0] sub_ln703_833_fu_2642_p2;
wire   [15:0] sub_ln703_834_fu_2646_p2;
wire   [15:0] sub_ln703_835_fu_2651_p2;
wire   [15:0] sub_ln703_836_fu_2655_p2;
wire   [15:0] sub_ln703_804_fu_2429_p2;
wire   [15:0] add_ln703_786_fu_3027_p2;
wire   [15:0] sub_ln703_837_fu_2660_p2;
wire   [15:0] sub_ln703_838_fu_2664_p2;
wire   [15:0] add_ln703_752_fu_2673_p2;
wire   [15:0] acc_1_V_fu_2678_p2;
wire   [15:0] acc_2_V_fu_2683_p2;
wire   [15:0] acc_3_V_fu_2688_p2;
wire   [15:0] acc_4_V_fu_2698_p2;
wire   [15:0] acc_5_V_fu_2703_p2;
wire   [15:0] acc_6_V_fu_2708_p2;
wire   [15:0] acc_7_V_fu_2713_p2;
wire   [15:0] acc_8_V_fu_2718_p2;
wire   [15:0] acc_9_V_fu_2723_p2;
wire   [15:0] acc_10_V_fu_2733_p2;
wire   [15:0] acc_11_V_fu_2738_p2;
wire   [15:0] acc_12_V_fu_2743_p2;
wire   [15:0] acc_13_V_fu_2748_p2;
wire   [15:0] acc_14_V_fu_2753_p2;
wire   [15:0] acc_15_V_fu_2758_p2;
wire   [15:0] acc_16_V_fu_2771_p2;
wire   [15:0] acc_17_V_fu_2777_p2;
wire   [15:0] acc_18_V_fu_2782_p2;
wire   [15:0] acc_19_V_fu_2787_p2;
wire   [15:0] acc_20_V_fu_2797_p2;
wire   [15:0] acc_21_V_fu_2802_p2;
wire   [15:0] acc_22_V_fu_2807_p2;
wire   [15:0] acc_23_V_fu_2812_p2;
wire   [15:0] acc_24_V_fu_2817_p2;
wire   [15:0] acc_25_V_fu_2822_p2;
wire   [15:0] acc_26_V_fu_2827_p2;
wire   [15:0] acc_27_V_fu_2832_p2;
wire   [15:0] acc_28_V_fu_2837_p2;
wire   [15:0] acc_29_V_fu_2842_p2;
wire   [15:0] acc_30_V_fu_2847_p2;
wire   [15:0] acc_31_V_fu_2852_p2;
wire   [15:0] acc_32_V_fu_2857_p2;
wire   [15:0] acc_33_V_fu_2862_p2;
wire   [15:0] acc_34_V_fu_2872_p2;
wire   [15:0] acc_35_V_fu_2877_p2;
wire   [15:0] acc_36_V_fu_2882_p2;
wire   [15:0] acc_37_V_fu_2887_p2;
wire   [15:0] acc_38_V_fu_2892_p2;
wire   [15:0] acc_39_V_fu_2897_p2;
wire   [15:0] acc_40_V_fu_2902_p2;
wire   [15:0] acc_41_V_fu_2907_p2;
wire   [15:0] acc_42_V_fu_2912_p2;
wire   [15:0] acc_43_V_fu_2917_p2;
wire   [15:0] acc_44_V_fu_2922_p2;
wire   [15:0] acc_45_V_fu_2927_p2;
wire   [15:0] acc_46_V_fu_2932_p2;
wire   [15:0] acc_47_V_fu_2942_p2;
wire   [15:0] acc_48_V_fu_2952_p2;
wire   [15:0] acc_49_V_fu_2962_p2;
wire   [15:0] acc_50_V_fu_2967_p2;
wire   [15:0] acc_51_V_fu_2972_p2;
wire   [15:0] acc_52_V_fu_2977_p2;
wire   [15:0] acc_53_V_fu_2982_p2;
wire   [15:0] acc_54_V_fu_2987_p2;
wire   [15:0] acc_55_V_fu_2997_p2;
wire   [15:0] acc_56_V_fu_3002_p2;
wire   [15:0] acc_57_V_fu_3007_p2;
wire   [15:0] acc_58_V_fu_3012_p2;
wire   [15:0] acc_59_V_fu_3017_p2;
wire   [15:0] acc_60_V_fu_3022_p2;
wire   [15:0] acc_61_V_fu_3031_p2;
wire   [15:0] acc_62_V_fu_3037_p2;
wire   [15:0] acc_63_V_fu_3042_p2;
reg    ap_ce_reg;
reg   [255:0] data_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;
reg   [15:0] ap_return_32_int_reg;
reg   [15:0] ap_return_33_int_reg;
reg   [15:0] ap_return_34_int_reg;
reg   [15:0] ap_return_35_int_reg;
reg   [15:0] ap_return_36_int_reg;
reg   [15:0] ap_return_37_int_reg;
reg   [15:0] ap_return_38_int_reg;
reg   [15:0] ap_return_39_int_reg;
reg   [15:0] ap_return_40_int_reg;
reg   [15:0] ap_return_41_int_reg;
reg   [15:0] ap_return_42_int_reg;
reg   [15:0] ap_return_43_int_reg;
reg   [15:0] ap_return_44_int_reg;
reg   [15:0] ap_return_45_int_reg;
reg   [15:0] ap_return_46_int_reg;
reg   [15:0] ap_return_47_int_reg;
reg   [15:0] ap_return_48_int_reg;
reg   [15:0] ap_return_49_int_reg;
reg   [15:0] ap_return_50_int_reg;
reg   [15:0] ap_return_51_int_reg;
reg   [15:0] ap_return_52_int_reg;
reg   [15:0] ap_return_53_int_reg;
reg   [15:0] ap_return_54_int_reg;
reg   [15:0] ap_return_55_int_reg;
reg   [15:0] ap_return_56_int_reg;
reg   [15:0] ap_return_57_int_reg;
reg   [15:0] ap_return_58_int_reg;
reg   [15:0] ap_return_59_int_reg;
reg   [15:0] ap_return_60_int_reg;
reg   [15:0] ap_return_61_int_reg;
reg   [15:0] ap_return_62_int_reg;
reg   [15:0] ap_return_63_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        add_ln703_538_reg_4067 <= add_ln703_538_fu_280_p2;
        add_ln703_538_reg_4067_pp0_iter4_reg <= add_ln703_538_reg_4067;
        add_ln703_539_reg_4035 <= add_ln703_539_fu_260_p2;
        add_ln703_539_reg_4035_pp0_iter2_reg <= add_ln703_539_reg_4035;
        add_ln703_539_reg_4035_pp0_iter3_reg <= add_ln703_539_reg_4035_pp0_iter2_reg;
        add_ln703_540_reg_4079 <= add_ln703_540_fu_288_p2;
        add_ln703_540_reg_4079_pp0_iter4_reg <= add_ln703_540_reg_4079;
        add_ln703_541_reg_4171 <= add_ln703_541_fu_348_p2;
        add_ln703_542_reg_4177 <= add_ln703_542_fu_352_p2;
        add_ln703_543_reg_4054 <= add_ln703_543_fu_272_p2;
        add_ln703_543_reg_4054_pp0_iter3_reg <= add_ln703_543_reg_4054;
        add_ln703_543_reg_4054_pp0_iter4_reg <= add_ln703_543_reg_4054_pp0_iter3_reg;
        add_ln703_544_reg_4116 <= add_ln703_544_fu_312_p2;
        add_ln703_544_reg_4116_pp0_iter5_reg <= add_ln703_544_reg_4116;
        add_ln703_545_reg_4183 <= add_ln703_545_fu_364_p2;
        add_ln703_547_reg_4128 <= add_ln703_547_fu_320_p2;
        add_ln703_548_reg_4188 <= add_ln703_548_fu_368_p2;
        add_ln703_549_reg_4103 <= add_ln703_549_fu_304_p2;
        add_ln703_549_reg_4103_pp0_iter4_reg <= add_ln703_549_reg_4103;
        add_ln703_549_reg_4103_pp0_iter5_reg <= add_ln703_549_reg_4103_pp0_iter4_reg;
        add_ln703_550_reg_4211 <= add_ln703_550_fu_384_p2;
        add_ln703_551_reg_4222 <= add_ln703_551_fu_393_p2;
        add_ln703_554_reg_4134 <= add_ln703_554_fu_324_p2;
        add_ln703_554_reg_4134_pp0_iter5_reg <= add_ln703_554_reg_4134;
        add_ln703_557_reg_4293 <= add_ln703_557_fu_488_p2;
        add_ln703_558_reg_4298 <= add_ln703_558_fu_498_p2;
        add_ln703_559_reg_4146 <= add_ln703_559_fu_332_p2;
        add_ln703_559_reg_4146_pp0_iter5_reg <= add_ln703_559_reg_4146;
        add_ln703_560_reg_4153 <= add_ln703_560_fu_336_p2;
        add_ln703_560_reg_4153_pp0_iter5_reg <= add_ln703_560_reg_4153;
        add_ln703_564_reg_4240 <= add_ln703_564_fu_406_p2;
        add_ln703_566_reg_4258 <= add_ln703_566_fu_418_p2;
        add_ln703_566_reg_4258_pp0_iter6_reg <= add_ln703_566_reg_4258;
        add_ln703_568_reg_4270 <= add_ln703_568_fu_426_p2;
        add_ln703_571_reg_4372 <= add_ln703_571_fu_657_p2;
        add_ln703_572_reg_4382 <= add_ln703_572_fu_670_p2;
        add_ln703_573_reg_4387 <= add_ln703_573_fu_675_p2;
        add_ln703_574_reg_4393 <= add_ln703_574_fu_679_p2;
        add_ln703_576_reg_4408 <= add_ln703_576_fu_702_p2;
        add_ln703_577_reg_4413 <= add_ln703_577_fu_707_p2;
        add_ln703_579_reg_4418 <= add_ln703_579_fu_716_p2;
        add_ln703_580_reg_4433 <= add_ln703_580_fu_730_p2;
        add_ln703_583_reg_4450 <= add_ln703_583_fu_754_p2;
        add_ln703_587_reg_4471 <= add_ln703_587_fu_786_p2;
        add_ln703_588_reg_4476 <= add_ln703_588_fu_792_p2;
        add_ln703_590_reg_4481 <= add_ln703_590_fu_801_p2;
        add_ln703_597_reg_4282 <= add_ln703_597_fu_434_p2;
        add_ln703_597_reg_4282_pp0_iter6_reg <= add_ln703_597_reg_4282;
        add_ln703_611_reg_4521 <= add_ln703_611_fu_887_p2;
        add_ln703_620_reg_4537 <= add_ln703_620_fu_891_p2;
        add_ln703_631_reg_4588 <= add_ln703_631_fu_1397_p2;
        add_ln703_634_reg_4593 <= add_ln703_634_fu_1416_p2;
        add_ln703_637_reg_4553 <= add_ln703_637_fu_906_p2;
        add_ln703_639_reg_4608 <= add_ln703_639_fu_1459_p2;
        add_ln703_642_reg_4628 <= add_ln703_642_fu_1505_p2;
        add_ln703_645_reg_4648 <= add_ln703_645_fu_1538_p2;
        add_ln703_646_reg_4658 <= add_ln703_646_fu_1553_p2;
        add_ln703_655_reg_4558 <= add_ln703_655_fu_910_p2;
        add_ln703_658_reg_4733 <= add_ln703_658_fu_1696_p2;
        add_ln703_659_reg_4568 <= add_ln703_659_fu_914_p2;
        add_ln703_661_reg_4744 <= add_ln703_661_fu_1710_p2;
        add_ln703_663_reg_4764 <= add_ln703_663_fu_1735_p2;
        add_ln703_667_reg_4784 <= add_ln703_667_fu_1767_p2;
        add_ln703_669_reg_4804 <= add_ln703_669_fu_1787_p2;
        add_ln703_670_reg_4819 <= add_ln703_670_fu_1802_p2;
        add_ln703_672_reg_4829 <= add_ln703_672_fu_1812_p2;
        add_ln703_674_reg_4839 <= add_ln703_674_fu_1822_p2;
        add_ln703_679_reg_4847 <= add_ln703_679_fu_1826_p2;
        add_ln703_687_reg_4857 <= add_ln703_687_fu_1847_p2;
        add_ln703_688_reg_4862 <= add_ln703_688_fu_1853_p2;
        add_ln703_692_reg_4573 <= add_ln703_692_fu_920_p2;
        add_ln703_692_reg_4573_pp0_iter7_reg <= add_ln703_692_reg_4573;
        add_ln703_707_reg_4867 <= add_ln703_707_fu_1877_p2;
        add_ln703_711_reg_4872 <= add_ln703_711_fu_1887_p2;
        add_ln703_716_reg_4877 <= add_ln703_716_fu_1902_p2;
        add_ln703_722_reg_4882 <= add_ln703_722_fu_1913_p2;
        add_ln703_724_reg_4887 <= add_ln703_724_fu_1923_p2;
        add_ln703_727_reg_4892 <= add_ln703_727_fu_1934_p2;
        add_ln703_729_reg_4897 <= add_ln703_729_fu_1945_p2;
        add_ln703_732_reg_4902 <= add_ln703_732_fu_1956_p2;
        add_ln703_737_reg_4907 <= add_ln703_737_fu_1962_p2;
        add_ln703_739_reg_4915 <= add_ln703_739_fu_1966_p2;
        add_ln703_751_reg_4920 <= add_ln703_751_fu_1971_p2;
        add_ln703_reg_4010 <= add_ln703_fu_242_p2;
        add_ln703_reg_4010_pp0_iter1_reg <= add_ln703_reg_4010;
        add_ln703_reg_4010_pp0_iter2_reg <= add_ln703_reg_4010_pp0_iter1_reg;
        mult_307_V_reg_3472 <= {{data_V_read_int_reg[79:64]}};
        mult_307_V_reg_3472_pp0_iter1_reg <= mult_307_V_reg_3472;
        mult_307_V_reg_3472_pp0_iter2_reg <= mult_307_V_reg_3472_pp0_iter1_reg;
        mult_307_V_reg_3472_pp0_iter3_reg <= mult_307_V_reg_3472_pp0_iter2_reg;
        mult_307_V_reg_3472_pp0_iter4_reg <= mult_307_V_reg_3472_pp0_iter3_reg;
        mult_307_V_reg_3472_pp0_iter5_reg <= mult_307_V_reg_3472_pp0_iter4_reg;
        mult_320_V_reg_3500 <= {{data_V_read_int_reg[95:80]}};
        mult_320_V_reg_3500_pp0_iter1_reg <= mult_320_V_reg_3500;
        mult_320_V_reg_3500_pp0_iter2_reg <= mult_320_V_reg_3500_pp0_iter1_reg;
        mult_320_V_reg_3500_pp0_iter3_reg <= mult_320_V_reg_3500_pp0_iter2_reg;
        mult_320_V_reg_3500_pp0_iter4_reg <= mult_320_V_reg_3500_pp0_iter3_reg;
        mult_320_V_reg_3500_pp0_iter5_reg <= mult_320_V_reg_3500_pp0_iter4_reg;
        mult_386_V_reg_3539 <= {{data_V_read_int_reg[111:96]}};
        mult_386_V_reg_3539_pp0_iter1_reg <= mult_386_V_reg_3539;
        mult_386_V_reg_3539_pp0_iter2_reg <= mult_386_V_reg_3539_pp0_iter1_reg;
        mult_386_V_reg_3539_pp0_iter3_reg <= mult_386_V_reg_3539_pp0_iter2_reg;
        mult_386_V_reg_3539_pp0_iter4_reg <= mult_386_V_reg_3539_pp0_iter3_reg;
        mult_386_V_reg_3539_pp0_iter5_reg <= mult_386_V_reg_3539_pp0_iter4_reg;
        mult_386_V_reg_3539_pp0_iter6_reg <= mult_386_V_reg_3539_pp0_iter5_reg;
        mult_449_V_reg_3582 <= {{data_V_read_int_reg[127:112]}};
        mult_449_V_reg_3582_pp0_iter1_reg <= mult_449_V_reg_3582;
        mult_449_V_reg_3582_pp0_iter2_reg <= mult_449_V_reg_3582_pp0_iter1_reg;
        mult_449_V_reg_3582_pp0_iter3_reg <= mult_449_V_reg_3582_pp0_iter2_reg;
        mult_449_V_reg_3582_pp0_iter4_reg <= mult_449_V_reg_3582_pp0_iter3_reg;
        mult_449_V_reg_3582_pp0_iter5_reg <= mult_449_V_reg_3582_pp0_iter4_reg;
        mult_449_V_reg_3582_pp0_iter6_reg <= mult_449_V_reg_3582_pp0_iter5_reg;
        mult_512_V_reg_3629 <= {{data_V_read_int_reg[143:128]}};
        mult_512_V_reg_3629_pp0_iter1_reg <= mult_512_V_reg_3629;
        mult_512_V_reg_3629_pp0_iter2_reg <= mult_512_V_reg_3629_pp0_iter1_reg;
        mult_512_V_reg_3629_pp0_iter3_reg <= mult_512_V_reg_3629_pp0_iter2_reg;
        mult_512_V_reg_3629_pp0_iter4_reg <= mult_512_V_reg_3629_pp0_iter3_reg;
        mult_512_V_reg_3629_pp0_iter5_reg <= mult_512_V_reg_3629_pp0_iter4_reg;
        mult_512_V_reg_3629_pp0_iter6_reg <= mult_512_V_reg_3629_pp0_iter5_reg;
        mult_576_V_reg_3674 <= {{data_V_read_int_reg[159:144]}};
        mult_576_V_reg_3674_pp0_iter1_reg <= mult_576_V_reg_3674;
        mult_576_V_reg_3674_pp0_iter2_reg <= mult_576_V_reg_3674_pp0_iter1_reg;
        mult_576_V_reg_3674_pp0_iter3_reg <= mult_576_V_reg_3674_pp0_iter2_reg;
        mult_576_V_reg_3674_pp0_iter4_reg <= mult_576_V_reg_3674_pp0_iter3_reg;
        mult_576_V_reg_3674_pp0_iter5_reg <= mult_576_V_reg_3674_pp0_iter4_reg;
        mult_576_V_reg_3674_pp0_iter6_reg <= mult_576_V_reg_3674_pp0_iter5_reg;
        mult_640_V_reg_3716 <= {{data_V_read_int_reg[175:160]}};
        mult_640_V_reg_3716_pp0_iter1_reg <= mult_640_V_reg_3716;
        mult_640_V_reg_3716_pp0_iter2_reg <= mult_640_V_reg_3716_pp0_iter1_reg;
        mult_640_V_reg_3716_pp0_iter3_reg <= mult_640_V_reg_3716_pp0_iter2_reg;
        mult_640_V_reg_3716_pp0_iter4_reg <= mult_640_V_reg_3716_pp0_iter3_reg;
        mult_640_V_reg_3716_pp0_iter5_reg <= mult_640_V_reg_3716_pp0_iter4_reg;
        mult_640_V_reg_3716_pp0_iter6_reg <= mult_640_V_reg_3716_pp0_iter5_reg;
        mult_704_V_reg_3765 <= {{data_V_read_int_reg[191:176]}};
        mult_704_V_reg_3765_pp0_iter1_reg <= mult_704_V_reg_3765;
        mult_704_V_reg_3765_pp0_iter2_reg <= mult_704_V_reg_3765_pp0_iter1_reg;
        mult_704_V_reg_3765_pp0_iter3_reg <= mult_704_V_reg_3765_pp0_iter2_reg;
        mult_704_V_reg_3765_pp0_iter4_reg <= mult_704_V_reg_3765_pp0_iter3_reg;
        mult_704_V_reg_3765_pp0_iter5_reg <= mult_704_V_reg_3765_pp0_iter4_reg;
        mult_704_V_reg_3765_pp0_iter6_reg <= mult_704_V_reg_3765_pp0_iter5_reg;
        mult_704_V_reg_3765_pp0_iter7_reg <= mult_704_V_reg_3765_pp0_iter6_reg;
        mult_770_V_reg_3814 <= {{data_V_read_int_reg[207:192]}};
        mult_770_V_reg_3814_pp0_iter1_reg <= mult_770_V_reg_3814;
        mult_770_V_reg_3814_pp0_iter2_reg <= mult_770_V_reg_3814_pp0_iter1_reg;
        mult_770_V_reg_3814_pp0_iter3_reg <= mult_770_V_reg_3814_pp0_iter2_reg;
        mult_770_V_reg_3814_pp0_iter4_reg <= mult_770_V_reg_3814_pp0_iter3_reg;
        mult_770_V_reg_3814_pp0_iter5_reg <= mult_770_V_reg_3814_pp0_iter4_reg;
        mult_770_V_reg_3814_pp0_iter6_reg <= mult_770_V_reg_3814_pp0_iter5_reg;
        mult_770_V_reg_3814_pp0_iter7_reg <= mult_770_V_reg_3814_pp0_iter6_reg;
        mult_832_V_reg_3861 <= {{data_V_read_int_reg[223:208]}};
        mult_832_V_reg_3861_pp0_iter1_reg <= mult_832_V_reg_3861;
        mult_832_V_reg_3861_pp0_iter2_reg <= mult_832_V_reg_3861_pp0_iter1_reg;
        mult_832_V_reg_3861_pp0_iter3_reg <= mult_832_V_reg_3861_pp0_iter2_reg;
        mult_832_V_reg_3861_pp0_iter4_reg <= mult_832_V_reg_3861_pp0_iter3_reg;
        mult_832_V_reg_3861_pp0_iter5_reg <= mult_832_V_reg_3861_pp0_iter4_reg;
        mult_832_V_reg_3861_pp0_iter6_reg <= mult_832_V_reg_3861_pp0_iter5_reg;
        mult_832_V_reg_3861_pp0_iter7_reg <= mult_832_V_reg_3861_pp0_iter6_reg;
        mult_896_V_reg_3909 <= {{data_V_read_int_reg[239:224]}};
        mult_896_V_reg_3909_pp0_iter1_reg <= mult_896_V_reg_3909;
        mult_896_V_reg_3909_pp0_iter2_reg <= mult_896_V_reg_3909_pp0_iter1_reg;
        mult_896_V_reg_3909_pp0_iter3_reg <= mult_896_V_reg_3909_pp0_iter2_reg;
        mult_896_V_reg_3909_pp0_iter4_reg <= mult_896_V_reg_3909_pp0_iter3_reg;
        mult_896_V_reg_3909_pp0_iter5_reg <= mult_896_V_reg_3909_pp0_iter4_reg;
        mult_896_V_reg_3909_pp0_iter6_reg <= mult_896_V_reg_3909_pp0_iter5_reg;
        mult_896_V_reg_3909_pp0_iter7_reg <= mult_896_V_reg_3909_pp0_iter6_reg;
        mult_960_V_reg_3958 <= {{data_V_read_int_reg[255:240]}};
        mult_960_V_reg_3958_pp0_iter1_reg <= mult_960_V_reg_3958;
        mult_960_V_reg_3958_pp0_iter2_reg <= mult_960_V_reg_3958_pp0_iter1_reg;
        mult_960_V_reg_3958_pp0_iter3_reg <= mult_960_V_reg_3958_pp0_iter2_reg;
        mult_960_V_reg_3958_pp0_iter4_reg <= mult_960_V_reg_3958_pp0_iter3_reg;
        mult_960_V_reg_3958_pp0_iter5_reg <= mult_960_V_reg_3958_pp0_iter4_reg;
        mult_960_V_reg_3958_pp0_iter6_reg <= mult_960_V_reg_3958_pp0_iter5_reg;
        mult_960_V_reg_3958_pp0_iter7_reg <= mult_960_V_reg_3958_pp0_iter6_reg;
        sub_ln703_531_reg_4023 <= sub_ln703_531_fu_252_p2;
        sub_ln703_531_reg_4023_pp0_iter2_reg <= sub_ln703_531_reg_4023;
        sub_ln703_532_reg_4061 <= sub_ln703_532_fu_276_p2;
        sub_ln703_532_reg_4061_pp0_iter4_reg <= sub_ln703_532_reg_4061;
        sub_ln703_533_reg_4042 <= sub_ln703_533_fu_264_p2;
        sub_ln703_533_reg_4042_pp0_iter3_reg <= sub_ln703_533_reg_4042;
        sub_ln703_533_reg_4042_pp0_iter4_reg <= sub_ln703_533_reg_4042_pp0_iter3_reg;
        sub_ln703_534_reg_4029 <= sub_ln703_534_fu_256_p2;
        sub_ln703_534_reg_4029_pp0_iter2_reg <= sub_ln703_534_reg_4029;
        sub_ln703_534_reg_4029_pp0_iter3_reg <= sub_ln703_534_reg_4029_pp0_iter2_reg;
        sub_ln703_534_reg_4029_pp0_iter4_reg <= sub_ln703_534_reg_4029_pp0_iter3_reg;
        sub_ln703_535_reg_4073 <= sub_ln703_535_fu_284_p2;
        sub_ln703_535_reg_4073_pp0_iter4_reg <= sub_ln703_535_reg_4073;
        sub_ln703_536_reg_4159 <= sub_ln703_536_fu_340_p2;
        sub_ln703_537_reg_4085 <= sub_ln703_537_fu_292_p2;
        sub_ln703_537_reg_4085_pp0_iter4_reg <= sub_ln703_537_reg_4085;
        sub_ln703_537_reg_4085_pp0_iter5_reg <= sub_ln703_537_reg_4085_pp0_iter4_reg;
        sub_ln703_538_reg_4048 <= sub_ln703_538_fu_268_p2;
        sub_ln703_538_reg_4048_pp0_iter3_reg <= sub_ln703_538_reg_4048;
        sub_ln703_538_reg_4048_pp0_iter4_reg <= sub_ln703_538_reg_4048_pp0_iter3_reg;
        sub_ln703_538_reg_4048_pp0_iter5_reg <= sub_ln703_538_reg_4048_pp0_iter4_reg;
        sub_ln703_539_reg_4165 <= sub_ln703_539_fu_344_p2;
        sub_ln703_540_reg_4110 <= sub_ln703_540_fu_308_p2;
        sub_ln703_540_reg_4110_pp0_iter5_reg <= sub_ln703_540_reg_4110;
        sub_ln703_543_reg_4091 <= sub_ln703_543_fu_296_p2;
        sub_ln703_543_reg_4091_pp0_iter4_reg <= sub_ln703_543_reg_4091;
        sub_ln703_544_reg_4122 <= sub_ln703_544_fu_316_p2;
        sub_ln703_544_reg_4122_pp0_iter5_reg <= sub_ln703_544_reg_4122;
        sub_ln703_545_reg_4097 <= sub_ln703_545_fu_300_p2;
        sub_ln703_545_reg_4097_pp0_iter4_reg <= sub_ln703_545_reg_4097;
        sub_ln703_545_reg_4097_pp0_iter5_reg <= sub_ln703_545_reg_4097_pp0_iter4_reg;
        sub_ln703_549_reg_4194 <= sub_ln703_549_fu_372_p2;
        sub_ln703_550_reg_4200 <= sub_ln703_550_fu_376_p2;
        sub_ln703_551_reg_4205 <= sub_ln703_551_fu_380_p2;
        sub_ln703_552_reg_4217 <= sub_ln703_552_fu_388_p2;
        sub_ln703_554_reg_4228 <= sub_ln703_554_fu_398_p2;
        sub_ln703_557_reg_4234 <= sub_ln703_557_fu_402_p2;
        sub_ln703_558_reg_4140 <= sub_ln703_558_fu_328_p2;
        sub_ln703_558_reg_4140_pp0_iter5_reg <= sub_ln703_558_reg_4140;
        sub_ln703_567_reg_4303 <= sub_ln703_567_fu_540_p2;
        sub_ln703_570_reg_4246 <= sub_ln703_570_fu_410_p2;
        sub_ln703_572_reg_4309 <= sub_ln703_572_fu_563_p2;
        sub_ln703_574_reg_4314 <= sub_ln703_574_fu_572_p2;
        sub_ln703_576_reg_4252 <= sub_ln703_576_fu_414_p2;
        sub_ln703_576_reg_4252_pp0_iter6_reg <= sub_ln703_576_reg_4252;
        sub_ln703_578_reg_4319 <= sub_ln703_578_fu_585_p2;
        sub_ln703_579_reg_4324 <= sub_ln703_579_fu_590_p2;
        sub_ln703_582_reg_4329 <= sub_ln703_582_fu_599_p2;
        sub_ln703_584_reg_4264 <= sub_ln703_584_fu_422_p2;
        sub_ln703_584_reg_4264_pp0_iter6_reg <= sub_ln703_584_reg_4264;
        sub_ln703_585_reg_4334 <= sub_ln703_585_fu_609_p2;
        sub_ln703_586_reg_4340 <= sub_ln703_586_fu_614_p2;
        sub_ln703_587_reg_4345 <= sub_ln703_587_fu_619_p2;
        sub_ln703_588_reg_4350 <= sub_ln703_588_fu_624_p2;
        sub_ln703_589_reg_4355 <= sub_ln703_589_fu_638_p2;
        sub_ln703_590_reg_4361 <= sub_ln703_590_fu_643_p2;
        sub_ln703_591_reg_4277 <= sub_ln703_591_fu_430_p2;
        sub_ln703_592_reg_4366 <= sub_ln703_592_fu_653_p2;
        sub_ln703_594_reg_4377 <= sub_ln703_594_fu_666_p2;
        sub_ln703_596_reg_4398 <= sub_ln703_596_fu_683_p2;
        sub_ln703_599_reg_4403 <= sub_ln703_599_fu_693_p2;
        sub_ln703_605_reg_4423 <= sub_ln703_605_fu_720_p2;
        sub_ln703_608_reg_4428 <= sub_ln703_608_fu_725_p2;
        sub_ln703_610_reg_4439 <= sub_ln703_610_fu_734_p2;
        sub_ln703_611_reg_4444 <= sub_ln703_611_fu_739_p2;
        sub_ln703_613_reg_4455 <= sub_ln703_613_fu_758_p2;
        sub_ln703_617_reg_4460 <= sub_ln703_617_fu_763_p2;
        sub_ln703_620_reg_4466 <= sub_ln703_620_fu_772_p2;
        sub_ln703_627_reg_4486 <= sub_ln703_627_fu_807_p2;
        sub_ln703_632_reg_4491 <= sub_ln703_632_fu_818_p2;
        sub_ln703_641_reg_4496 <= sub_ln703_641_fu_838_p2;
        sub_ln703_645_reg_4501 <= sub_ln703_645_fu_843_p2;
        sub_ln703_660_reg_4506 <= sub_ln703_660_fu_872_p2;
        sub_ln703_661_reg_4511 <= sub_ln703_661_fu_877_p2;
        sub_ln703_662_reg_4516 <= sub_ln703_662_fu_882_p2;
        sub_ln703_671_reg_4543 <= sub_ln703_671_fu_896_p2;
        sub_ln703_676_reg_4548 <= sub_ln703_676_fu_901_p2;
        sub_ln703_692_reg_4598 <= sub_ln703_692_fu_1433_p2;
        sub_ln703_693_reg_4603 <= sub_ln703_693_fu_1438_p2;
        sub_ln703_695_reg_4613 <= sub_ln703_695_fu_1464_p2;
        sub_ln703_699_reg_4618 <= sub_ln703_699_fu_1495_p2;
        sub_ln703_700_reg_4623 <= sub_ln703_700_fu_1500_p2;
        sub_ln703_701_reg_4633 <= sub_ln703_701_fu_1509_p2;
        sub_ln703_702_reg_4638 <= sub_ln703_702_fu_1514_p2;
        sub_ln703_704_reg_4643 <= sub_ln703_704_fu_1524_p2;
        sub_ln703_706_reg_4653 <= sub_ln703_706_fu_1548_p2;
        sub_ln703_707_reg_4663 <= sub_ln703_707_fu_1559_p2;
        sub_ln703_708_reg_4668 <= sub_ln703_708_fu_1564_p2;
        sub_ln703_709_reg_4673 <= sub_ln703_709_fu_1569_p2;
        sub_ln703_710_reg_4678 <= sub_ln703_710_fu_1606_p2;
        sub_ln703_711_reg_4683 <= sub_ln703_711_fu_1611_p2;
        sub_ln703_712_reg_4688 <= sub_ln703_712_fu_1616_p2;
        sub_ln703_714_reg_4693 <= sub_ln703_714_fu_1626_p2;
        sub_ln703_715_reg_4698 <= sub_ln703_715_fu_1631_p2;
        sub_ln703_716_reg_4703 <= sub_ln703_716_fu_1636_p2;
        sub_ln703_718_reg_4708 <= sub_ln703_718_fu_1646_p2;
        sub_ln703_720_reg_4713 <= sub_ln703_720_fu_1676_p2;
        sub_ln703_722_reg_4718 <= sub_ln703_722_fu_1681_p2;
        sub_ln703_724_reg_4723 <= sub_ln703_724_fu_1686_p2;
        sub_ln703_725_reg_4728 <= sub_ln703_725_fu_1691_p2;
        sub_ln703_727_reg_4738 <= sub_ln703_727_fu_1701_p2;
        sub_ln703_729_reg_4749 <= sub_ln703_729_fu_1715_p2;
        sub_ln703_730_reg_4754 <= sub_ln703_730_fu_1720_p2;
        sub_ln703_731_reg_4759 <= sub_ln703_731_fu_1725_p2;
        sub_ln703_732_reg_4769 <= sub_ln703_732_fu_1741_p2;
        sub_ln703_738_reg_4774 <= sub_ln703_738_fu_1757_p2;
        sub_ln703_742_reg_4779 <= sub_ln703_742_fu_1762_p2;
        sub_ln703_743_reg_4789 <= sub_ln703_743_fu_1772_p2;
        sub_ln703_744_reg_4794 <= sub_ln703_744_fu_1777_p2;
        sub_ln703_745_reg_4799 <= sub_ln703_745_fu_1782_p2;
        sub_ln703_748_reg_4809 <= sub_ln703_748_fu_1792_p2;
        sub_ln703_751_reg_4814 <= sub_ln703_751_fu_1797_p2;
        sub_ln703_752_reg_4824 <= sub_ln703_752_fu_1807_p2;
        sub_ln703_753_reg_4834 <= sub_ln703_753_fu_1817_p2;
        sub_ln703_765_reg_4852 <= sub_ln703_765_fu_1832_p2;
        sub_ln703_reg_4017 <= sub_ln703_fu_248_p2;
        sub_ln703_reg_4017_pp0_iter2_reg <= sub_ln703_reg_4017;
        tmp_2_reg_3437 <= {{data_V_read_int_reg[31:16]}};
        tmp_3_reg_3443 <= {{data_V_read_int_reg[47:32]}};
        tmp_3_reg_3443_pp0_iter1_reg <= tmp_3_reg_3443;
        tmp_3_reg_3443_pp0_iter2_reg <= tmp_3_reg_3443_pp0_iter1_reg;
        tmp_4_reg_3454 <= {{data_V_read_int_reg[63:48]}};
        tmp_4_reg_3454_pp0_iter1_reg <= tmp_4_reg_3454;
        tmp_4_reg_3454_pp0_iter2_reg <= tmp_4_reg_3454_pp0_iter1_reg;
        tmp_4_reg_3454_pp0_iter3_reg <= tmp_4_reg_3454_pp0_iter2_reg;
        tmp_4_reg_3454_pp0_iter4_reg <= tmp_4_reg_3454_pp0_iter3_reg;
        trunc_ln203_reg_3431 <= trunc_ln203_fu_88_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_752_fu_2673_p2;
        ap_return_10_int_reg <= acc_10_V_fu_2733_p2;
        ap_return_11_int_reg <= acc_11_V_fu_2738_p2;
        ap_return_12_int_reg <= acc_12_V_fu_2743_p2;
        ap_return_13_int_reg <= acc_13_V_fu_2748_p2;
        ap_return_14_int_reg <= acc_14_V_fu_2753_p2;
        ap_return_15_int_reg <= acc_15_V_fu_2758_p2;
        ap_return_16_int_reg <= acc_16_V_fu_2771_p2;
        ap_return_17_int_reg <= acc_17_V_fu_2777_p2;
        ap_return_18_int_reg <= acc_18_V_fu_2782_p2;
        ap_return_19_int_reg <= acc_19_V_fu_2787_p2;
        ap_return_1_int_reg <= acc_1_V_fu_2678_p2;
        ap_return_20_int_reg <= acc_20_V_fu_2797_p2;
        ap_return_21_int_reg <= acc_21_V_fu_2802_p2;
        ap_return_22_int_reg <= acc_22_V_fu_2807_p2;
        ap_return_23_int_reg <= acc_23_V_fu_2812_p2;
        ap_return_24_int_reg <= acc_24_V_fu_2817_p2;
        ap_return_25_int_reg <= acc_25_V_fu_2822_p2;
        ap_return_26_int_reg <= acc_26_V_fu_2827_p2;
        ap_return_27_int_reg <= acc_27_V_fu_2832_p2;
        ap_return_28_int_reg <= acc_28_V_fu_2837_p2;
        ap_return_29_int_reg <= acc_29_V_fu_2842_p2;
        ap_return_2_int_reg <= acc_2_V_fu_2683_p2;
        ap_return_30_int_reg <= acc_30_V_fu_2847_p2;
        ap_return_31_int_reg <= acc_31_V_fu_2852_p2;
        ap_return_32_int_reg <= acc_32_V_fu_2857_p2;
        ap_return_33_int_reg <= acc_33_V_fu_2862_p2;
        ap_return_34_int_reg <= acc_34_V_fu_2872_p2;
        ap_return_35_int_reg <= acc_35_V_fu_2877_p2;
        ap_return_36_int_reg <= acc_36_V_fu_2882_p2;
        ap_return_37_int_reg <= acc_37_V_fu_2887_p2;
        ap_return_38_int_reg <= acc_38_V_fu_2892_p2;
        ap_return_39_int_reg <= acc_39_V_fu_2897_p2;
        ap_return_3_int_reg <= acc_3_V_fu_2688_p2;
        ap_return_40_int_reg <= acc_40_V_fu_2902_p2;
        ap_return_41_int_reg <= acc_41_V_fu_2907_p2;
        ap_return_42_int_reg <= acc_42_V_fu_2912_p2;
        ap_return_43_int_reg <= acc_43_V_fu_2917_p2;
        ap_return_44_int_reg <= acc_44_V_fu_2922_p2;
        ap_return_45_int_reg <= acc_45_V_fu_2927_p2;
        ap_return_46_int_reg <= acc_46_V_fu_2932_p2;
        ap_return_47_int_reg <= acc_47_V_fu_2942_p2;
        ap_return_48_int_reg <= acc_48_V_fu_2952_p2;
        ap_return_49_int_reg <= acc_49_V_fu_2962_p2;
        ap_return_4_int_reg <= acc_4_V_fu_2698_p2;
        ap_return_50_int_reg <= acc_50_V_fu_2967_p2;
        ap_return_51_int_reg <= acc_51_V_fu_2972_p2;
        ap_return_52_int_reg <= acc_52_V_fu_2977_p2;
        ap_return_53_int_reg <= acc_53_V_fu_2982_p2;
        ap_return_54_int_reg <= acc_54_V_fu_2987_p2;
        ap_return_55_int_reg <= acc_55_V_fu_2997_p2;
        ap_return_56_int_reg <= acc_56_V_fu_3002_p2;
        ap_return_57_int_reg <= acc_57_V_fu_3007_p2;
        ap_return_58_int_reg <= acc_58_V_fu_3012_p2;
        ap_return_59_int_reg <= acc_59_V_fu_3017_p2;
        ap_return_5_int_reg <= acc_5_V_fu_2703_p2;
        ap_return_60_int_reg <= acc_60_V_fu_3022_p2;
        ap_return_61_int_reg <= acc_61_V_fu_3031_p2;
        ap_return_62_int_reg <= acc_62_V_fu_3037_p2;
        ap_return_63_int_reg <= acc_63_V_fu_3042_p2;
        ap_return_6_int_reg <= acc_6_V_fu_2708_p2;
        ap_return_7_int_reg <= acc_7_V_fu_2713_p2;
        ap_return_8_int_reg <= acc_8_V_fu_2718_p2;
        ap_return_9_int_reg <= acc_9_V_fu_2723_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_V_read_int_reg <= data_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_752_fu_2673_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_2678_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = acc_10_V_fu_2733_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = acc_11_V_fu_2738_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = acc_12_V_fu_2743_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = acc_13_V_fu_2748_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = acc_14_V_fu_2753_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = acc_15_V_fu_2758_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = acc_16_V_fu_2771_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = acc_17_V_fu_2777_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = acc_18_V_fu_2782_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = acc_19_V_fu_2787_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_2683_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = acc_20_V_fu_2797_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = acc_21_V_fu_2802_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = acc_22_V_fu_2807_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = acc_23_V_fu_2812_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = acc_24_V_fu_2817_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = acc_25_V_fu_2822_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = acc_26_V_fu_2827_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = acc_27_V_fu_2832_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = acc_28_V_fu_2837_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = acc_29_V_fu_2842_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_2688_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = acc_30_V_fu_2847_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = acc_31_V_fu_2852_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_32 = ap_return_32_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_32 = acc_32_V_fu_2857_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_33 = ap_return_33_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_33 = acc_33_V_fu_2862_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_34 = ap_return_34_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_34 = acc_34_V_fu_2872_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_35 = ap_return_35_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_35 = acc_35_V_fu_2877_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_36 = ap_return_36_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_36 = acc_36_V_fu_2882_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_37 = ap_return_37_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_37 = acc_37_V_fu_2887_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_38 = ap_return_38_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_38 = acc_38_V_fu_2892_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_39 = ap_return_39_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_39 = acc_39_V_fu_2897_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_2698_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_40 = ap_return_40_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_40 = acc_40_V_fu_2902_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_41 = ap_return_41_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_41 = acc_41_V_fu_2907_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_42 = ap_return_42_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_42 = acc_42_V_fu_2912_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_43 = ap_return_43_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_43 = acc_43_V_fu_2917_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_44 = ap_return_44_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_44 = acc_44_V_fu_2922_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_45 = ap_return_45_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_45 = acc_45_V_fu_2927_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_46 = ap_return_46_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_46 = acc_46_V_fu_2932_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_47 = ap_return_47_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_47 = acc_47_V_fu_2942_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_48 = ap_return_48_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_48 = acc_48_V_fu_2952_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_49 = ap_return_49_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_49 = acc_49_V_fu_2962_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = acc_5_V_fu_2703_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_50 = ap_return_50_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_50 = acc_50_V_fu_2967_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_51 = ap_return_51_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_51 = acc_51_V_fu_2972_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_52 = ap_return_52_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_52 = acc_52_V_fu_2977_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_53 = ap_return_53_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_53 = acc_53_V_fu_2982_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_54 = ap_return_54_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_54 = acc_54_V_fu_2987_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_55 = ap_return_55_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_55 = acc_55_V_fu_2997_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_56 = ap_return_56_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_56 = acc_56_V_fu_3002_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_57 = ap_return_57_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_57 = acc_57_V_fu_3007_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_58 = ap_return_58_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_58 = acc_58_V_fu_3012_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_59 = ap_return_59_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_59 = acc_59_V_fu_3017_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = acc_6_V_fu_2708_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_60 = ap_return_60_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_60 = acc_60_V_fu_3022_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_61 = ap_return_61_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_61 = acc_61_V_fu_3031_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_62 = ap_return_62_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_62 = acc_62_V_fu_3037_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_63 = ap_return_63_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_63 = acc_63_V_fu_3042_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = acc_7_V_fu_2713_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = acc_8_V_fu_2718_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = acc_9_V_fu_2723_p2;
    end
end

assign acc_10_V_fu_2733_p2 = (add_ln703_758_fu_2728_p2 + add_ln703_751_reg_4920);

assign acc_11_V_fu_2738_p2 = (sub_ln703_811_fu_2474_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_12_V_fu_2743_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_812_fu_2479_p2);

assign acc_13_V_fu_2748_p2 = (add_ln703_735_fu_2484_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_14_V_fu_2753_p2 = (sub_ln703_813_fu_2489_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_15_V_fu_2758_p2 = (sub_ln703_814_fu_2494_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_16_V_fu_2771_p2 = (add_ln703_761_fu_2763_p2 + add_ln703_762_fu_2767_p2);

assign acc_17_V_fu_2777_p2 = (sub_ln703_815_fu_2499_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_18_V_fu_2782_p2 = (add_ln703_736_fu_2504_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_19_V_fu_2787_p2 = (sub_ln703_790_fu_2299_p2 + add_ln703_751_reg_4920);

assign acc_1_V_fu_2678_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_805_fu_2439_p2);

assign acc_20_V_fu_2797_p2 = (add_ln703_765_fu_2792_p2 + add_ln703_751_reg_4920);

assign acc_21_V_fu_2802_p2 = (sub_ln703_816_fu_2509_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_22_V_fu_2807_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_817_fu_2514_p2);

assign acc_23_V_fu_2812_p2 = (sub_ln703_818_fu_2519_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_24_V_fu_2817_p2 = (sub_ln703_819_fu_2524_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_25_V_fu_2822_p2 = (sub_ln703_791_fu_2318_p2 + add_ln703_751_reg_4920);

assign acc_26_V_fu_2827_p2 = (add_ln703_738_fu_2528_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_27_V_fu_2832_p2 = (add_ln703_741_fu_2536_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_28_V_fu_2837_p2 = (sub_ln703_820_fu_2541_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_29_V_fu_2842_p2 = (sub_ln703_821_fu_2546_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_2_V_fu_2683_p2 = (sub_ln703_806_fu_2444_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_30_V_fu_2847_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_822_fu_2550_p2);

assign acc_31_V_fu_2852_p2 = (sub_ln703_823_fu_2555_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_32_V_fu_2857_p2 = (sub_ln703_824_fu_2560_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_33_V_fu_2862_p2 = (sub_ln703_825_fu_2564_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_34_V_fu_2872_p2 = (add_ln703_770_fu_2867_p2 + add_ln703_751_reg_4920);

assign acc_35_V_fu_2877_p2 = (add_ln703_742_fu_2569_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_36_V_fu_2882_p2 = (sub_ln703_793_fu_2356_p2 + add_ln703_751_reg_4920);

assign acc_37_V_fu_2887_p2 = (sub_ln703_826_fu_2574_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_38_V_fu_2892_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_827_fu_2579_p2);

assign acc_39_V_fu_2897_p2 = (add_ln703_743_fu_2583_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_3_V_fu_2688_p2 = (sub_ln703_807_fu_2449_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_40_V_fu_2902_p2 = (sub_ln703_828_fu_2588_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_41_V_fu_2907_p2 = (sub_ln703_829_fu_2593_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_42_V_fu_2912_p2 = (sub_ln703_830_fu_2598_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_43_V_fu_2917_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_831_fu_2602_p2);

assign acc_44_V_fu_2922_p2 = (sub_ln703_797_fu_2385_p2 + add_ln703_751_reg_4920);

assign acc_45_V_fu_2927_p2 = (sub_ln703_832_fu_2607_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_46_V_fu_2932_p2 = (add_ln703_744_fu_2612_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_47_V_fu_2942_p2 = (add_ln703_776_fu_2937_p2 + add_ln703_751_reg_4920);

assign acc_48_V_fu_2952_p2 = (add_ln703_778_fu_2947_p2 + add_ln703_751_reg_4920);

assign acc_49_V_fu_2962_p2 = (add_ln703_780_fu_2957_p2 + add_ln703_751_reg_4920);

assign acc_4_V_fu_2698_p2 = (add_ln703_754_fu_2693_p2 + add_ln703_751_reg_4920);

assign acc_50_V_fu_2967_p2 = (add_ln703_745_fu_2617_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_51_V_fu_2972_p2 = (add_ln703_746_fu_2622_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_52_V_fu_2977_p2 = (add_ln703_747_fu_2627_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_53_V_fu_2982_p2 = (add_ln703_748_fu_2632_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_54_V_fu_2987_p2 = (add_ln703_749_fu_2637_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_55_V_fu_2997_p2 = (add_ln703_782_fu_2992_p2 + add_ln703_751_reg_4920);

assign acc_56_V_fu_3002_p2 = (sub_ln703_833_fu_2642_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_57_V_fu_3007_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_834_fu_2646_p2);

assign acc_58_V_fu_3012_p2 = (sub_ln703_835_fu_2651_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_59_V_fu_3017_p2 = (sub_ln703_836_fu_2655_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_5_V_fu_2703_p2 = (sub_ln703_808_fu_2454_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_60_V_fu_3022_p2 = (sub_ln703_804_fu_2429_p2 + add_ln703_751_reg_4920);

assign acc_61_V_fu_3031_p2 = (add_ln703_786_fu_3027_p2 + add_ln703_762_fu_2767_p2);

assign acc_62_V_fu_3037_p2 = (sub_ln703_837_fu_2660_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_63_V_fu_3042_p2 = (sub_ln703_838_fu_2664_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_6_V_fu_2708_p2 = (sub_ln703_809_fu_2459_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_7_V_fu_2713_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_810_fu_2464_p2);

assign acc_8_V_fu_2718_p2 = (sub_ln703_785_fu_2254_p2 + add_ln703_751_reg_4920);

assign acc_9_V_fu_2723_p2 = (add_ln703_734_fu_2469_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign add_ln703_538_fu_280_p2 = (tmp_3_reg_3443_pp0_iter2_reg + sub_ln703_reg_4017_pp0_iter2_reg);

assign add_ln703_539_fu_260_p2 = (tmp_3_reg_3443 + add_ln703_reg_4010);

assign add_ln703_540_fu_288_p2 = (tmp_3_reg_3443_pp0_iter2_reg + sub_ln703_531_reg_4023_pp0_iter2_reg);

assign add_ln703_541_fu_348_p2 = (tmp_4_reg_3454_pp0_iter4_reg + sub_ln703_535_reg_4073_pp0_iter4_reg);

assign add_ln703_542_fu_352_p2 = (tmp_4_reg_3454_pp0_iter4_reg + sub_ln703_534_reg_4029_pp0_iter4_reg);

assign add_ln703_543_fu_272_p2 = (tmp_4_reg_3454_pp0_iter1_reg + add_ln703_539_reg_4035);

assign add_ln703_544_fu_312_p2 = (tmp_4_reg_3454_pp0_iter3_reg + sub_ln703_532_reg_4061);

assign add_ln703_545_fu_364_p2 = (tmp_4_reg_3454_pp0_iter4_reg + sub_ln703_533_reg_4042_pp0_iter4_reg);

assign add_ln703_546_fu_438_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_536_reg_4159);

assign add_ln703_547_fu_320_p2 = (mult_307_V_reg_3472_pp0_iter3_reg + tmp_4_reg_3454_pp0_iter3_reg);

assign add_ln703_548_fu_368_p2 = (add_ln703_538_reg_4067_pp0_iter4_reg + add_ln703_547_reg_4128);

assign add_ln703_549_fu_304_p2 = (mult_307_V_reg_3472_pp0_iter2_reg + add_ln703_543_reg_4054);

assign add_ln703_550_fu_384_p2 = (add_ln703_540_reg_4079_pp0_iter4_reg + add_ln703_547_reg_4128);

assign add_ln703_551_fu_393_p2 = (mult_307_V_reg_3472_pp0_iter4_reg + sub_ln703_542_fu_360_p2);

assign add_ln703_552_fu_454_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + add_ln703_542_reg_4177);

assign add_ln703_553_fu_458_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_539_reg_4165);

assign add_ln703_554_fu_324_p2 = (mult_307_V_reg_3472_pp0_iter3_reg + sub_ln703_543_reg_4091);

assign add_ln703_555_fu_466_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_538_reg_4048_pp0_iter5_reg);

assign add_ln703_556_fu_478_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_546_fu_438_p2);

assign add_ln703_557_fu_488_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_547_fu_446_p2);

assign add_ln703_558_fu_498_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_548_reg_4188);

assign add_ln703_559_fu_332_p2 = (mult_320_V_reg_3500_pp0_iter3_reg + add_ln703_549_reg_4103);

assign add_ln703_560_fu_336_p2 = (mult_320_V_reg_3500_pp0_iter3_reg + mult_307_V_reg_3472_pp0_iter3_reg);

assign add_ln703_561_fu_510_p2 = (add_ln703_541_reg_4171 + add_ln703_560_reg_4153_pp0_iter5_reg);

assign add_ln703_562_fu_522_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_552_reg_4217);

assign add_ln703_563_fu_526_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_551_reg_4222);

assign add_ln703_564_fu_406_p2 = (add_ln703_544_reg_4116 + add_ln703_560_reg_4153);

assign add_ln703_565_fu_554_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_544_reg_4122_pp0_iter5_reg);

assign add_ln703_566_fu_418_p2 = (mult_386_V_reg_3539_pp0_iter4_reg + sub_ln703_558_reg_4140);

assign add_ln703_567_fu_629_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_537_reg_4085_pp0_iter5_reg);

assign add_ln703_568_fu_426_p2 = (mult_386_V_reg_3539_pp0_iter4_reg + mult_320_V_reg_3500_pp0_iter4_reg);

assign add_ln703_569_fu_633_p2 = (add_ln703_567_fu_629_p2 + add_ln703_568_reg_4270);

assign add_ln703_570_fu_648_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_566_fu_535_p2);

assign add_ln703_571_fu_657_p2 = (sub_ln703_554_reg_4228 + add_ln703_568_reg_4270);

assign add_ln703_572_fu_670_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_569_fu_549_p2);

assign add_ln703_573_fu_675_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + add_ln703_559_reg_4146_pp0_iter5_reg);

assign add_ln703_574_fu_679_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_570_reg_4246);

assign add_ln703_575_fu_698_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + add_ln703_564_reg_4240);

assign add_ln703_576_fu_702_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_575_fu_577_p2);

assign add_ln703_577_fu_707_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_577_fu_581_p2);

assign add_ln703_578_fu_944_p2 = (mult_386_V_reg_3539_pp0_iter6_reg + add_ln703_558_reg_4298);

assign add_ln703_579_fu_716_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_576_reg_4252);

assign add_ln703_580_fu_730_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + sub_ln703_584_reg_4264);

assign add_ln703_581_fu_744_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + mult_386_V_reg_3539_pp0_iter5_reg);

assign add_ln703_582_fu_748_p2 = (sub_ln703_564_fu_518_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_583_fu_754_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + add_ln703_566_reg_4258);

assign add_ln703_584_fu_985_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_592_reg_4366);

assign add_ln703_585_fu_777_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_540_reg_4110_pp0_iter5_reg);

assign add_ln703_586_fu_781_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_581_fu_744_p2);

assign add_ln703_587_fu_786_p2 = (add_ln703_585_fu_777_p2 + add_ln703_586_fu_781_p2);

assign add_ln703_588_fu_792_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + sub_ln703_597_fu_688_p2);

assign add_ln703_589_fu_797_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_545_reg_4097_pp0_iter5_reg);

assign add_ln703_590_fu_801_p2 = (add_ln703_589_fu_797_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_591_fu_1027_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + add_ln703_573_reg_4387);

assign add_ln703_592_fu_1031_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_589_reg_4355);

assign add_ln703_593_fu_812_p2 = (sub_ln703_568_fu_545_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_594_fu_823_p2 = (sub_ln703_557_reg_4234 + add_ln703_581_fu_744_p2);

assign add_ln703_595_fu_828_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_550_reg_4211);

assign add_ln703_596_fu_832_p2 = (add_ln703_595_fu_828_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_597_fu_434_p2 = (mult_512_V_reg_3629_pp0_iter4_reg + mult_449_V_reg_3582_pp0_iter4_reg);

assign add_ln703_598_fu_1052_p2 = (sub_ln703_579_reg_4324 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_599_fu_1073_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_609_fu_965_p2);

assign add_ln703_600_fu_848_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_554_reg_4134_pp0_iter5_reg);

assign add_ln703_601_fu_852_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + add_ln703_597_reg_4282);

assign add_ln703_602_fu_856_p2 = (add_ln703_600_fu_848_p2 + add_ln703_601_fu_852_p2);

assign add_ln703_603_fu_1132_p2 = (sub_ln703_596_reg_4398 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_604_fu_1140_p2 = (sub_ln703_598_fu_932_p2 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_605_fu_862_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_549_reg_4194);

assign add_ln703_606_fu_866_p2 = (add_ln703_605_fu_862_p2 + add_ln703_601_fu_852_p2);

assign add_ln703_607_fu_1163_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_611_reg_4444);

assign add_ln703_608_fu_1176_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_631_fu_1039_p2);

assign add_ln703_609_fu_1181_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_632_reg_4491);

assign add_ln703_610_fu_1185_p2 = (sub_ln703_586_reg_4340 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_611_fu_887_p2 = (mult_576_V_reg_3674_pp0_iter5_reg + mult_512_V_reg_3629_pp0_iter5_reg);

assign add_ln703_612_fu_1194_p2 = (sub_ln703_604_fu_952_p2 + add_ln703_611_reg_4521);

assign add_ln703_613_fu_1209_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_638_fu_1069_p2);

assign add_ln703_614_fu_1219_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_639_fu_1078_p2);

assign add_ln703_615_fu_1228_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_643_fu_1091_p2);

assign add_ln703_616_fu_1238_p2 = (sub_ln703_615_fu_977_p2 + add_ln703_611_reg_4521);

assign add_ln703_617_fu_1243_p2 = (sub_ln703_616_fu_981_p2 + add_ln703_611_reg_4521);

assign add_ln703_618_fu_1248_p2 = (add_ln703_580_reg_4433 + add_ln703_611_reg_4521);

assign add_ln703_619_fu_1252_p2 = (sub_ln703_617_reg_4460 + add_ln703_611_reg_4521);

assign add_ln703_620_fu_891_p2 = (mult_576_V_reg_3674_pp0_iter5_reg + sub_ln703_645_fu_843_p2);

assign add_ln703_621_fu_1256_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_646_fu_1099_p2);

assign add_ln703_622_fu_1271_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_648_fu_1108_p2);

assign add_ln703_623_fu_1276_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_649_fu_1113_p2);

assign add_ln703_624_fu_1286_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_652_fu_1127_p2);

assign add_ln703_625_fu_1311_p2 = (sub_ln703_629_fu_1022_p2 + add_ln703_611_reg_4521);

assign add_ln703_626_fu_1321_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_587_reg_4345);

assign add_ln703_627_fu_1325_p2 = (add_ln703_626_fu_1321_p2 + add_ln703_611_reg_4521);

assign add_ln703_628_fu_1350_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_601_fu_940_p2);

assign add_ln703_629_fu_1355_p2 = (add_ln703_628_fu_1350_p2 + add_ln703_611_reg_4521);

assign add_ln703_630_fu_1387_p2 = (sub_ln703_634_fu_1048_p2 + add_ln703_611_reg_4521);

assign add_ln703_631_fu_1397_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + add_ln703_612_fu_1194_p2);

assign add_ln703_632_fu_1407_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_606_fu_956_p2);

assign add_ln703_633_fu_1412_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + mult_576_V_reg_3674_pp0_iter6_reg);

assign add_ln703_634_fu_1416_p2 = (add_ln703_632_fu_1407_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_635_fu_1422_p2 = (sub_ln703_636_fu_1060_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_636_fu_1448_p2 = (sub_ln703_640_fu_1082_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_637_fu_906_p2 = (sub_ln703_551_reg_4205 + add_ln703_568_reg_4270);

assign add_ln703_638_fu_1454_p2 = (add_ln703_597_reg_4282_pp0_iter6_reg + add_ln703_633_fu_1412_p2);

assign add_ln703_639_fu_1459_p2 = (add_ln703_637_reg_4553 + add_ln703_638_fu_1454_p2);

assign add_ln703_640_fu_1469_p2 = (sub_ln703_642_fu_1086_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_641_fu_1480_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_668_fu_1233_p2);

assign add_ln703_642_fu_1505_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + add_ln703_620_reg_4537);

assign add_ln703_643_fu_1529_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_585_reg_4334);

assign add_ln703_644_fu_1533_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + add_ln703_633_fu_1412_p2);

assign add_ln703_645_fu_1538_p2 = (add_ln703_643_fu_1529_p2 + add_ln703_644_fu_1533_p2);

assign add_ln703_646_fu_1553_p2 = (sub_ln703_650_fu_1118_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_647_fu_1574_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_674_fu_1296_p2);

assign add_ln703_648_fu_1579_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_626_fu_1014_p2);

assign add_ln703_649_fu_1584_p2 = (add_ln703_648_fu_1579_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_650_fu_1590_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_677_fu_1306_p2);

assign add_ln703_651_fu_1595_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_628_fu_1018_p2);

assign add_ln703_652_fu_1600_p2 = (add_ln703_651_fu_1595_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_653_fu_1651_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_687_fu_1378_p2);

assign add_ln703_654_fu_1661_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_603_fu_948_p2);

assign add_ln703_655_fu_910_p2 = (mult_704_V_reg_3765_pp0_iter5_reg + mult_640_V_reg_3716_pp0_iter5_reg);

assign add_ln703_656_fu_1666_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + add_ln703_655_reg_4558);

assign add_ln703_657_fu_1670_p2 = (add_ln703_654_fu_1661_p2 + add_ln703_656_fu_1666_p2);

assign add_ln703_658_fu_1696_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + sub_ln703_694_fu_1443_p2);

assign add_ln703_659_fu_914_p2 = (sub_ln703_563_fu_514_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_660_fu_1706_p2 = (add_ln703_611_reg_4521 + add_ln703_655_reg_4558);

assign add_ln703_661_fu_1710_p2 = (add_ln703_659_reg_4568 + add_ln703_660_fu_1706_p2);

assign add_ln703_662_fu_1730_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_614_fu_973_p2);

assign add_ln703_663_fu_1735_p2 = (add_ln703_662_fu_1730_p2 + add_ln703_656_fu_1666_p2);

assign add_ln703_664_fu_1991_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_699_reg_4618);

assign add_ln703_665_fu_1746_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_619_fu_989_p2);

assign add_ln703_666_fu_1751_p2 = (add_ln703_665_fu_1746_p2 + add_ln703_656_fu_1666_p2);

assign add_ln703_667_fu_1767_p2 = (sub_ln703_675_fu_1301_p2 + add_ln703_655_reg_4558);

assign add_ln703_668_fu_2035_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_712_reg_4688);

assign add_ln703_669_fu_1787_p2 = (sub_ln703_680_fu_1335_p2 + add_ln703_655_reg_4558);

assign add_ln703_670_fu_1802_p2 = (sub_ln703_685_fu_1370_p2 + add_ln703_655_reg_4558);

assign add_ln703_671_fu_2047_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_718_reg_4708);

assign add_ln703_672_fu_1812_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + sub_ln703_719_fu_1656_p2);

assign add_ln703_673_fu_2068_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_725_reg_4728);

assign add_ln703_674_fu_1822_p2 = (mult_770_V_reg_3814_pp0_iter6_reg + mult_704_V_reg_3765_pp0_iter6_reg);

assign add_ln703_675_fu_2072_p2 = (sub_ln703_692_reg_4598 + add_ln703_674_reg_4839);

assign add_ln703_676_fu_2093_p2 = (sub_ln703_695_reg_4613 + add_ln703_674_reg_4839);

assign add_ln703_677_fu_2101_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_730_reg_4754);

assign add_ln703_678_fu_2109_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_732_reg_4769);

assign add_ln703_679_fu_1826_p2 = (sub_ln703_698_fu_1490_p2 + add_ln703_674_fu_1822_p2);

assign add_ln703_680_fu_2118_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_736_fu_2007_p2);

assign add_ln703_681_fu_2132_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_727_reg_4738);

assign add_ln703_682_fu_2136_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_740_fu_2019_p2);

assign add_ln703_683_fu_2146_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_742_reg_4779);

assign add_ln703_684_fu_2154_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_743_reg_4789);

assign add_ln703_685_fu_1837_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_654_fu_1145_p2);

assign add_ln703_686_fu_1842_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + add_ln703_674_fu_1822_p2);

assign add_ln703_687_fu_1847_p2 = (add_ln703_685_fu_1837_p2 + add_ln703_686_fu_1842_p2);

assign add_ln703_688_fu_1853_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_679_fu_1330_p2);

assign add_ln703_689_fu_2181_p2 = (add_ln703_688_reg_4862 + add_ln703_674_reg_4839);

assign add_ln703_690_fu_2189_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_748_reg_4809);

assign add_ln703_691_fu_2193_p2 = (sub_ln703_714_reg_4693 + add_ln703_674_reg_4839);

assign add_ln703_692_fu_920_p2 = (mult_832_V_reg_3861_pp0_iter5_reg + mult_770_V_reg_3814_pp0_iter5_reg);

assign add_ln703_693_fu_2229_p2 = (sub_ln703_721_fu_1975_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_694_fu_2234_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_755_fu_2055_p2);

assign add_ln703_695_fu_2239_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_757_fu_2064_p2);

assign add_ln703_696_fu_2264_p2 = (sub_ln703_728_fu_1987_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_697_fu_2269_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_761_fu_2089_p2);

assign add_ln703_698_fu_2279_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_762_fu_2097_p2);

assign add_ln703_699_fu_2289_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_763_fu_2105_p2);

assign add_ln703_700_fu_2303_p2 = (sub_ln703_733_fu_1995_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_701_fu_2308_p2 = (sub_ln703_734_fu_1999_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_702_fu_2313_p2 = (sub_ln703_735_fu_2003_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_703_fu_1858_p2 = (mult_386_V_reg_3539_pp0_iter6_reg + sub_ln703_567_reg_4303);

assign add_ln703_704_fu_1862_p2 = (add_ln703_703_fu_1858_p2 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_705_fu_1867_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + add_ln703_692_reg_4573);

assign add_ln703_706_fu_1871_p2 = (add_ln703_633_fu_1412_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_707_fu_1877_p2 = (add_ln703_704_fu_1862_p2 + add_ln703_706_fu_1871_p2);

assign add_ln703_708_fu_2323_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_704_reg_4643);

assign add_ln703_709_fu_2327_p2 = (add_ln703_708_fu_2323_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_710_fu_1883_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_671_reg_4543);

assign add_ln703_711_fu_1887_p2 = (add_ln703_710_fu_1883_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_712_fu_2332_p2 = (sub_ln703_737_fu_2011_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_713_fu_2337_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_766_fu_2123_p2);

assign add_ln703_714_fu_1893_p2 = (sub_ln703_622_fu_997_p2 + add_ln703_611_reg_4521);

assign add_ln703_715_fu_1898_p2 = (add_ln703_655_reg_4558 + add_ln703_692_reg_4573);

assign add_ln703_716_fu_1902_p2 = (add_ln703_714_fu_1893_p2 + add_ln703_715_fu_1898_p2);

assign add_ln703_717_fu_2342_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_706_reg_4653);

assign add_ln703_718_fu_2346_p2 = (add_ln703_717_fu_2342_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_719_fu_2361_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_708_reg_4668);

assign add_ln703_720_fu_2365_p2 = (add_ln703_719_fu_2361_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_721_fu_1908_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_673_fu_1291_p2);

assign add_ln703_722_fu_1913_p2 = (add_ln703_721_fu_1908_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_723_fu_1919_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_676_reg_4548);

assign add_ln703_724_fu_1923_p2 = (add_ln703_723_fu_1919_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_725_fu_2389_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_770_fu_2158_p2);

assign add_ln703_726_fu_1929_p2 = (sub_ln703_660_reg_4506 + add_ln703_633_fu_1412_p2);

assign add_ln703_727_fu_1934_p2 = (add_ln703_726_fu_1929_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_728_fu_1940_p2 = (sub_ln703_633_fu_1043_p2 + add_ln703_611_reg_4521);

assign add_ln703_729_fu_1945_p2 = (add_ln703_728_fu_1940_p2 + add_ln703_715_fu_1898_p2);

assign add_ln703_730_fu_2424_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_779_fu_2211_p2);

assign add_ln703_731_fu_1951_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_688_fu_1382_p2);

assign add_ln703_732_fu_1956_p2 = (add_ln703_731_fu_1951_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_733_fu_2434_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_781_fu_2220_p2);

assign add_ln703_734_fu_2469_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_786_fu_2259_p2);

assign add_ln703_735_fu_2484_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_787_fu_2274_p2);

assign add_ln703_736_fu_2504_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_789_fu_2294_p2);

assign add_ln703_737_fu_1962_p2 = (mult_896_V_reg_3909_pp0_iter6_reg + mult_832_V_reg_3861_pp0_iter6_reg);

assign add_ln703_738_fu_2528_p2 = (sub_ln703_765_reg_4852 + add_ln703_737_reg_4907);

assign add_ln703_739_fu_1966_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + sub_ln703_703_fu_1519_p2);

assign add_ln703_740_fu_2532_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + add_ln703_737_reg_4907);

assign add_ln703_741_fu_2536_p2 = (add_ln703_739_reg_4915 + add_ln703_740_fu_2532_p2);

assign add_ln703_742_fu_2569_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_792_fu_2351_p2);

assign add_ln703_743_fu_2583_p2 = (sub_ln703_768_fu_2141_p2 + add_ln703_737_reg_4907);

assign add_ln703_744_fu_2612_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_798_fu_2394_p2);

assign add_ln703_745_fu_2617_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_799_fu_2399_p2);

assign add_ln703_746_fu_2622_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_800_fu_2404_p2);

assign add_ln703_747_fu_2627_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_801_fu_2409_p2);

assign add_ln703_748_fu_2632_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_802_fu_2414_p2);

assign add_ln703_749_fu_2637_p2 = (sub_ln703_776_fu_2197_p2 + add_ln703_737_reg_4907);

assign add_ln703_750_fu_2669_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_753_reg_4834);

assign add_ln703_751_fu_1971_p2 = (mult_960_V_reg_3958_pp0_iter6_reg + mult_896_V_reg_3909_pp0_iter6_reg);

assign add_ln703_752_fu_2673_p2 = (add_ln703_750_fu_2669_p2 + add_ln703_751_reg_4920);

assign add_ln703_754_fu_2693_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_756_fu_2059_p2);

assign add_ln703_758_fu_2728_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_760_fu_2085_p2);

assign add_ln703_761_fu_2763_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_731_reg_4759);

assign add_ln703_762_fu_2767_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + add_ln703_751_reg_4920);

assign add_ln703_765_fu_2792_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_764_fu_2113_p2);

assign add_ln703_770_fu_2867_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_767_fu_2127_p2);

assign add_ln703_776_fu_2937_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_772_fu_2166_p2);

assign add_ln703_778_fu_2947_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_773_fu_2171_p2);

assign add_ln703_780_fu_2957_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_774_fu_2176_p2);

assign add_ln703_782_fu_2992_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_777_fu_2202_p2);

assign add_ln703_786_fu_3027_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_752_reg_4824);

assign add_ln703_fu_242_p2 = (tmp_2_fu_92_p4 + trunc_ln203_fu_88_p1);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign sub_ln703_531_fu_252_p2 = (tmp_2_reg_3437 - trunc_ln203_reg_3431);

assign sub_ln703_532_fu_276_p2 = (sub_ln703_reg_4017_pp0_iter2_reg - tmp_3_reg_3443_pp0_iter2_reg);

assign sub_ln703_533_fu_264_p2 = (sub_ln703_531_reg_4023 - tmp_3_reg_3443_pp0_iter1_reg);

assign sub_ln703_534_fu_256_p2 = (add_ln703_reg_4010 - tmp_3_reg_3443);

assign sub_ln703_535_fu_284_p2 = (tmp_3_reg_3443_pp0_iter2_reg - add_ln703_reg_4010_pp0_iter2_reg);

assign sub_ln703_536_fu_340_p2 = (sub_ln703_532_reg_4061_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_537_fu_292_p2 = (sub_ln703_533_reg_4042 - tmp_4_reg_3454_pp0_iter2_reg);

assign sub_ln703_538_fu_268_p2 = (sub_ln703_534_reg_4029 - tmp_4_reg_3454_pp0_iter1_reg);

assign sub_ln703_539_fu_344_p2 = (add_ln703_538_reg_4067_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_540_fu_308_p2 = (tmp_4_reg_3454_pp0_iter3_reg - add_ln703_539_reg_4035_pp0_iter3_reg);

assign sub_ln703_541_fu_356_p2 = (add_ln703_540_reg_4079_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_542_fu_360_p2 = (sub_ln703_535_reg_4073_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_543_fu_296_p2 = (add_ln703_539_reg_4035_pp0_iter2_reg - tmp_4_reg_3454_pp0_iter2_reg);

assign sub_ln703_544_fu_316_p2 = (sub_ln703_537_reg_4085 - mult_307_V_reg_3472_pp0_iter3_reg);

assign sub_ln703_545_fu_300_p2 = (sub_ln703_538_reg_4048 - mult_307_V_reg_3472_pp0_iter2_reg);

assign sub_ln703_546_fu_442_p2 = (sub_ln703_539_reg_4165 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_547_fu_446_p2 = (add_ln703_541_reg_4171 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_548_fu_450_p2 = (add_ln703_542_reg_4177 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_549_fu_372_p2 = (add_ln703_543_reg_4054_pp0_iter4_reg - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_550_fu_376_p2 = (mult_307_V_reg_3472_pp0_iter4_reg - add_ln703_543_reg_4054_pp0_iter4_reg);

assign sub_ln703_551_fu_380_p2 = (sub_ln703_540_reg_4110 - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_552_fu_388_p2 = (sub_ln703_541_fu_356_p2 - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_553_fu_462_p2 = (add_ln703_544_reg_4116_pp0_iter5_reg - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_554_fu_398_p2 = (sub_ln703_543_reg_4091_pp0_iter4_reg - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_555_fu_470_p2 = (sub_ln703_536_reg_4159 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_556_fu_474_p2 = (add_ln703_545_reg_4183 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_557_fu_402_p2 = (sub_ln703_544_reg_4122 - mult_320_V_reg_3500_pp0_iter4_reg);

assign sub_ln703_558_fu_328_p2 = (sub_ln703_545_reg_4097 - mult_320_V_reg_3500_pp0_iter3_reg);

assign sub_ln703_559_fu_483_p2 = (sub_ln703_546_fu_442_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_560_fu_493_p2 = (sub_ln703_548_fu_450_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_561_fu_502_p2 = (sub_ln703_549_reg_4194 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_562_fu_506_p2 = (sub_ln703_550_reg_4200 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_563_fu_514_p2 = (add_ln703_550_reg_4211 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_564_fu_518_p2 = (mult_320_V_reg_3500_pp0_iter5_reg - add_ln703_549_reg_4103_pp0_iter5_reg);

assign sub_ln703_565_fu_530_p2 = (add_ln703_552_fu_454_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_566_fu_535_p2 = (add_ln703_553_fu_458_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_567_fu_540_p2 = (sub_ln703_553_fu_462_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_568_fu_545_p2 = (sub_ln703_551_reg_4205 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_569_fu_549_p2 = (add_ln703_546_fu_438_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_570_fu_410_p2 = (add_ln703_554_reg_4134 - mult_320_V_reg_3500_pp0_iter4_reg);

assign sub_ln703_571_fu_558_p2 = (add_ln703_555_fu_466_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_572_fu_563_p2 = (sub_ln703_554_reg_4228 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_573_fu_567_p2 = (sub_ln703_555_fu_470_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_574_fu_572_p2 = (sub_ln703_556_fu_474_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_575_fu_577_p2 = (add_ln703_548_reg_4188 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_576_fu_414_p2 = (add_ln703_549_reg_4103_pp0_iter4_reg - mult_320_V_reg_3500_pp0_iter4_reg);

assign sub_ln703_577_fu_581_p2 = (add_ln703_551_reg_4222 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_578_fu_585_p2 = (add_ln703_556_fu_478_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_579_fu_590_p2 = (sub_ln703_557_reg_4234 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_580_fu_594_p2 = (sub_ln703_559_fu_483_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_581_fu_924_p2 = (add_ln703_557_reg_4293 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_582_fu_599_p2 = (sub_ln703_560_fu_493_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_583_fu_604_p2 = (add_ln703_558_fu_498_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_584_fu_422_p2 = (add_ln703_559_reg_4146 - mult_386_V_reg_3539_pp0_iter4_reg);

assign sub_ln703_585_fu_609_p2 = (sub_ln703_561_fu_502_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_586_fu_614_p2 = (sub_ln703_562_fu_506_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_587_fu_619_p2 = (add_ln703_561_fu_510_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_588_fu_624_p2 = (add_ln703_562_fu_522_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_589_fu_638_p2 = (add_ln703_563_fu_526_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_590_fu_643_p2 = (sub_ln703_565_fu_530_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_591_fu_430_p2 = (mult_386_V_reg_3539_pp0_iter4_reg - add_ln703_559_reg_4146);

assign sub_ln703_592_fu_653_p2 = (sub_ln703_558_reg_4140_pp0_iter5_reg - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_593_fu_661_p2 = (sub_ln703_568_fu_545_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_594_fu_666_p2 = (add_ln703_564_reg_4240 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_595_fu_928_p2 = (sub_ln703_567_reg_4303 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_596_fu_683_p2 = (add_ln703_565_fu_554_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_597_fu_688_p2 = (sub_ln703_571_fu_558_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_598_fu_932_p2 = (sub_ln703_572_reg_4309 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_599_fu_693_p2 = (sub_ln703_573_fu_567_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_600_fu_936_p2 = (sub_ln703_574_reg_4314 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_601_fu_940_p2 = (sub_ln703_576_reg_4252_pp0_iter6_reg - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_602_fu_712_p2 = (sub_ln703_570_reg_4246 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_603_fu_948_p2 = (sub_ln703_578_reg_4319 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_604_fu_952_p2 = (add_ln703_566_reg_4258_pp0_iter6_reg - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_605_fu_720_p2 = (sub_ln703_580_fu_594_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_606_fu_956_p2 = (sub_ln703_581_fu_924_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_607_fu_961_p2 = (sub_ln703_582_reg_4329 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_608_fu_725_p2 = (sub_ln703_583_fu_604_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_609_fu_965_p2 = (sub_ln703_585_reg_4334 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_610_fu_734_p2 = (sub_ln703_586_fu_614_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_611_fu_739_p2 = (sub_ln703_587_fu_619_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_612_fu_969_p2 = (sub_ln703_588_reg_4350 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_613_fu_758_p2 = (add_ln703_569_fu_633_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_614_fu_973_p2 = (sub_ln703_589_reg_4355 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_615_fu_977_p2 = (sub_ln703_590_reg_4361 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_616_fu_981_p2 = (sub_ln703_584_reg_4264_pp0_iter6_reg - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_617_fu_763_p2 = (add_ln703_570_fu_648_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_618_fu_768_p2 = (sub_ln703_591_reg_4277 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_619_fu_989_p2 = (add_ln703_571_reg_4372 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_620_fu_772_p2 = (sub_ln703_593_fu_661_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_621_fu_993_p2 = (sub_ln703_594_reg_4377 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_622_fu_997_p2 = (sub_ln703_595_fu_928_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_623_fu_1002_p2 = (add_ln703_572_reg_4382 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_624_fu_1006_p2 = (add_ln703_573_reg_4387 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_625_fu_1010_p2 = (add_ln703_574_reg_4393 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_626_fu_1014_p2 = (sub_ln703_599_reg_4403 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_627_fu_807_p2 = (add_ln703_575_fu_698_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_628_fu_1018_p2 = (sub_ln703_592_reg_4366 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_629_fu_1022_p2 = (sub_ln703_600_fu_936_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_630_fu_1035_p2 = (add_ln703_576_reg_4408 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_631_fu_1039_p2 = (add_ln703_577_reg_4413 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_632_fu_818_p2 = (sub_ln703_602_fu_712_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_633_fu_1043_p2 = (add_ln703_578_fu_944_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_634_fu_1048_p2 = (add_ln703_579_reg_4418 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_635_fu_1056_p2 = (sub_ln703_605_reg_4423 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_636_fu_1060_p2 = (sub_ln703_607_fu_961_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_637_fu_1065_p2 = (sub_ln703_608_reg_4428 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_638_fu_1069_p2 = (add_ln703_580_reg_4433 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_639_fu_1078_p2 = (sub_ln703_610_reg_4439 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_640_fu_1082_p2 = (sub_ln703_611_reg_4444 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_641_fu_838_p2 = (add_ln703_582_fu_748_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_642_fu_1086_p2 = (sub_ln703_612_fu_969_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_643_fu_1091_p2 = (add_ln703_583_reg_4450 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_644_fu_1095_p2 = (sub_ln703_613_reg_4455 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_645_fu_843_p2 = (sub_ln703_618_fu_768_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_646_fu_1099_p2 = (add_ln703_584_fu_985_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_647_fu_1104_p2 = (sub_ln703_620_reg_4466 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_648_fu_1108_p2 = (sub_ln703_621_fu_993_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_649_fu_1113_p2 = (sub_ln703_623_fu_1002_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_650_fu_1118_p2 = (add_ln703_587_reg_4471 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_651_fu_1122_p2 = (sub_ln703_624_fu_1006_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_652_fu_1127_p2 = (sub_ln703_625_fu_1010_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_653_fu_1136_p2 = (add_ln703_588_reg_4476 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_654_fu_1145_p2 = (add_ln703_590_reg_4481 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_655_fu_1149_p2 = (sub_ln703_627_reg_4486 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_656_fu_1153_p2 = (add_ln703_591_fu_1027_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_657_fu_1158_p2 = (add_ln703_592_fu_1031_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_658_fu_1167_p2 = (sub_ln703_617_reg_4460 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_659_fu_1171_p2 = (sub_ln703_630_fu_1035_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_660_fu_872_p2 = (add_ln703_593_fu_812_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_661_fu_877_p2 = (add_ln703_594_fu_823_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_662_fu_882_p2 = (add_ln703_596_fu_832_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_663_fu_1189_p2 = (add_ln703_598_fu_1052_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_664_fu_1199_p2 = (sub_ln703_635_fu_1056_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_665_fu_1204_p2 = (sub_ln703_637_fu_1065_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_666_fu_1214_p2 = (add_ln703_599_fu_1073_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_667_fu_1224_p2 = (sub_ln703_641_reg_4496 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_668_fu_1233_p2 = (sub_ln703_644_fu_1095_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_669_fu_1261_p2 = (sub_ln703_636_fu_1060_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_670_fu_1266_p2 = (sub_ln703_647_fu_1104_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_671_fu_896_p2 = (add_ln703_602_fu_856_p2 - mult_576_V_reg_3674_pp0_iter5_reg);

assign sub_ln703_672_fu_1281_p2 = (sub_ln703_651_fu_1122_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_673_fu_1291_p2 = (add_ln703_603_fu_1132_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_674_fu_1296_p2 = (sub_ln703_653_fu_1136_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_675_fu_1301_p2 = (add_ln703_604_fu_1140_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_676_fu_901_p2 = (add_ln703_606_fu_866_p2 - mult_576_V_reg_3674_pp0_iter5_reg);

assign sub_ln703_677_fu_1306_p2 = (sub_ln703_655_fu_1149_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_678_fu_1316_p2 = (sub_ln703_656_fu_1153_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_679_fu_1330_p2 = (sub_ln703_657_fu_1158_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_680_fu_1335_p2 = (add_ln703_607_fu_1163_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_681_fu_1340_p2 = (sub_ln703_658_fu_1167_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_682_fu_1345_p2 = (sub_ln703_659_fu_1171_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_683_fu_1360_p2 = (add_ln703_608_fu_1176_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_684_fu_1365_p2 = (add_ln703_609_fu_1181_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_685_fu_1370_p2 = (sub_ln703_661_reg_4511 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_686_fu_1374_p2 = (sub_ln703_662_reg_4516 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_687_fu_1378_p2 = (sub_ln703_645_reg_4501 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_688_fu_1382_p2 = (add_ln703_610_fu_1185_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_689_fu_1392_p2 = (sub_ln703_663_fu_1189_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_690_fu_1402_p2 = (sub_ln703_664_fu_1199_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_691_fu_1428_p2 = (sub_ln703_665_fu_1204_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_692_fu_1433_p2 = (add_ln703_613_fu_1209_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_693_fu_1438_p2 = (sub_ln703_666_fu_1214_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_694_fu_1443_p2 = (add_ln703_614_fu_1219_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_695_fu_1464_p2 = (sub_ln703_667_fu_1224_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_696_fu_1475_p2 = (add_ln703_615_fu_1228_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_697_fu_1485_p2 = (add_ln703_616_fu_1238_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_698_fu_1490_p2 = (add_ln703_617_fu_1243_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_699_fu_1495_p2 = (add_ln703_618_fu_1248_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_700_fu_1500_p2 = (add_ln703_619_fu_1252_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_701_fu_1509_p2 = (add_ln703_621_fu_1256_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_702_fu_1514_p2 = (sub_ln703_669_fu_1261_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_703_fu_1519_p2 = (sub_ln703_670_fu_1266_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_704_fu_1524_p2 = (add_ln703_622_fu_1271_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_705_fu_1544_p2 = (add_ln703_620_reg_4537 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_706_fu_1548_p2 = (add_ln703_623_fu_1276_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_707_fu_1559_p2 = (sub_ln703_672_fu_1281_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_708_fu_1564_p2 = (add_ln703_624_fu_1286_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_709_fu_1569_p2 = (add_ln703_612_fu_1194_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_710_fu_1606_p2 = (add_ln703_625_fu_1311_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_711_fu_1611_p2 = (sub_ln703_678_fu_1316_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_712_fu_1616_p2 = (add_ln703_627_fu_1325_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_713_fu_1621_p2 = (sub_ln703_681_fu_1340_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_714_fu_1626_p2 = (sub_ln703_682_fu_1345_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_715_fu_1631_p2 = (add_ln703_629_fu_1355_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_716_fu_1636_p2 = (sub_ln703_683_fu_1360_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_717_fu_1641_p2 = (sub_ln703_684_fu_1365_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_718_fu_1646_p2 = (sub_ln703_686_fu_1374_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_719_fu_1656_p2 = (add_ln703_630_fu_1387_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_720_fu_1676_p2 = (sub_ln703_689_fu_1392_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_721_fu_1975_p2 = (add_ln703_631_reg_4588 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_722_fu_1681_p2 = (sub_ln703_690_fu_1402_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_723_fu_1979_p2 = (add_ln703_634_reg_4593 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_724_fu_1686_p2 = (add_ln703_635_fu_1422_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_725_fu_1691_p2 = (sub_ln703_691_fu_1428_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_726_fu_1983_p2 = (sub_ln703_693_reg_4603 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_727_fu_1701_p2 = (add_ln703_636_fu_1448_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_728_fu_1987_p2 = (add_ln703_639_reg_4608 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_729_fu_1715_p2 = (add_ln703_640_fu_1469_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_730_fu_1720_p2 = (sub_ln703_696_fu_1475_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_731_fu_1725_p2 = (add_ln703_641_fu_1480_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_732_fu_1741_p2 = (sub_ln703_697_fu_1485_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_733_fu_1995_p2 = (sub_ln703_700_reg_4623 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_734_fu_1999_p2 = (add_ln703_642_reg_4628 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_735_fu_2003_p2 = (sub_ln703_701_reg_4633 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_736_fu_2007_p2 = (sub_ln703_702_reg_4638 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_737_fu_2011_p2 = (add_ln703_645_reg_4648 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_738_fu_1757_p2 = (sub_ln703_705_fu_1544_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_739_fu_2015_p2 = (add_ln703_646_reg_4658 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_740_fu_2019_p2 = (sub_ln703_707_reg_4663 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_741_fu_2023_p2 = (sub_ln703_709_reg_4673 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_742_fu_1762_p2 = (add_ln703_647_fu_1574_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_743_fu_1772_p2 = (add_ln703_649_fu_1584_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_744_fu_1777_p2 = (add_ln703_650_fu_1590_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_745_fu_1782_p2 = (add_ln703_652_fu_1600_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_746_fu_2027_p2 = (sub_ln703_710_reg_4678 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_747_fu_2031_p2 = (sub_ln703_711_reg_4683 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_748_fu_1792_p2 = (sub_ln703_713_fu_1621_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_749_fu_2039_p2 = (sub_ln703_715_reg_4698 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_750_fu_2043_p2 = (sub_ln703_716_reg_4703 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_751_fu_1797_p2 = (sub_ln703_717_fu_1641_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_752_fu_1807_p2 = (add_ln703_653_fu_1651_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_753_fu_1817_p2 = (add_ln703_657_fu_1670_p2 - mult_770_V_reg_3814_pp0_iter6_reg);

assign sub_ln703_754_fu_2051_p2 = (sub_ln703_720_reg_4713 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_755_fu_2055_p2 = (sub_ln703_722_reg_4718 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_756_fu_2059_p2 = (sub_ln703_723_fu_1979_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_757_fu_2064_p2 = (sub_ln703_724_reg_4723 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_758_fu_2076_p2 = (sub_ln703_726_fu_1983_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_759_fu_2081_p2 = (add_ln703_658_reg_4733 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_760_fu_2085_p2 = (sub_ln703_727_reg_4738 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_761_fu_2089_p2 = (add_ln703_661_reg_4744 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_762_fu_2097_p2 = (sub_ln703_729_reg_4749 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_763_fu_2105_p2 = (add_ln703_663_reg_4764 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_764_fu_2113_p2 = (add_ln703_664_fu_1991_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_765_fu_1832_p2 = (add_ln703_666_fu_1751_p2 - mult_770_V_reg_3814_pp0_iter6_reg);

assign sub_ln703_766_fu_2123_p2 = (sub_ln703_738_reg_4774 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_767_fu_2127_p2 = (sub_ln703_739_fu_2015_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_768_fu_2141_p2 = (sub_ln703_741_fu_2023_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_769_fu_2150_p2 = (add_ln703_667_reg_4784 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_770_fu_2158_p2 = (sub_ln703_744_reg_4794 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_771_fu_2162_p2 = (sub_ln703_745_reg_4799 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_772_fu_2166_p2 = (sub_ln703_746_fu_2027_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_773_fu_2171_p2 = (sub_ln703_747_fu_2031_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_774_fu_2176_p2 = (add_ln703_668_fu_2035_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_775_fu_2185_p2 = (add_ln703_669_reg_4804 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_776_fu_2197_p2 = (sub_ln703_749_fu_2039_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_777_fu_2202_p2 = (sub_ln703_750_fu_2043_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_778_fu_2207_p2 = (sub_ln703_751_reg_4814 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_779_fu_2211_p2 = (add_ln703_670_reg_4819 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_780_fu_2215_p2 = (add_ln703_671_fu_2047_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_781_fu_2220_p2 = (add_ln703_672_reg_4829 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_782_fu_2224_p2 = (sub_ln703_754_fu_2051_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_783_fu_2244_p2 = (add_ln703_673_fu_2068_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_784_fu_2249_p2 = (add_ln703_675_fu_2072_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_785_fu_2254_p2 = (sub_ln703_758_fu_2076_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_786_fu_2259_p2 = (sub_ln703_759_fu_2081_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_787_fu_2274_p2 = (add_ln703_676_fu_2093_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_788_fu_2284_p2 = (add_ln703_677_fu_2101_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_789_fu_2294_p2 = (add_ln703_678_fu_2109_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_790_fu_2299_p2 = (add_ln703_679_reg_4847 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_791_fu_2318_p2 = (add_ln703_680_fu_2118_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_792_fu_2351_p2 = (add_ln703_681_fu_2132_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_793_fu_2356_p2 = (add_ln703_682_fu_2136_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_794_fu_2370_p2 = (add_ln703_683_fu_2146_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_795_fu_2375_p2 = (sub_ln703_769_fu_2150_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_796_fu_2380_p2 = (add_ln703_684_fu_2154_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_797_fu_2385_p2 = (add_ln703_687_reg_4857 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_798_fu_2394_p2 = (sub_ln703_771_fu_2162_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_799_fu_2399_p2 = (add_ln703_689_fu_2181_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_800_fu_2404_p2 = (sub_ln703_775_fu_2185_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_801_fu_2409_p2 = (add_ln703_690_fu_2189_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_802_fu_2414_p2 = (add_ln703_691_fu_2193_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_803_fu_2419_p2 = (sub_ln703_778_fu_2207_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_804_fu_2429_p2 = (sub_ln703_780_fu_2215_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_805_fu_2439_p2 = (sub_ln703_782_fu_2224_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_806_fu_2444_p2 = (add_ln703_693_fu_2229_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_807_fu_2449_p2 = (add_ln703_694_fu_2234_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_808_fu_2454_p2 = (add_ln703_695_fu_2239_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_809_fu_2459_p2 = (sub_ln703_783_fu_2244_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_810_fu_2464_p2 = (sub_ln703_784_fu_2249_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_811_fu_2474_p2 = (add_ln703_696_fu_2264_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_812_fu_2479_p2 = (add_ln703_697_fu_2269_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_813_fu_2489_p2 = (add_ln703_698_fu_2279_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_814_fu_2494_p2 = (sub_ln703_788_fu_2284_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_815_fu_2499_p2 = (add_ln703_699_fu_2289_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_816_fu_2509_p2 = (add_ln703_700_fu_2303_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_817_fu_2514_p2 = (add_ln703_701_fu_2308_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_818_fu_2519_p2 = (add_ln703_702_fu_2313_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_819_fu_2524_p2 = (add_ln703_707_reg_4867 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_820_fu_2541_p2 = (add_ln703_709_fu_2327_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_821_fu_2546_p2 = (add_ln703_711_reg_4872 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_822_fu_2550_p2 = (add_ln703_712_fu_2332_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_823_fu_2555_p2 = (add_ln703_713_fu_2337_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_824_fu_2560_p2 = (add_ln703_716_reg_4877 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_825_fu_2564_p2 = (add_ln703_718_fu_2346_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_826_fu_2574_p2 = (add_ln703_720_fu_2365_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_827_fu_2579_p2 = (add_ln703_722_reg_4882 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_828_fu_2588_p2 = (sub_ln703_794_fu_2370_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_829_fu_2593_p2 = (sub_ln703_795_fu_2375_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_830_fu_2598_p2 = (add_ln703_724_reg_4887 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_831_fu_2602_p2 = (sub_ln703_796_fu_2380_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_832_fu_2607_p2 = (add_ln703_725_fu_2389_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_833_fu_2642_p2 = (add_ln703_727_reg_4892 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_834_fu_2646_p2 = (sub_ln703_803_fu_2419_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_835_fu_2651_p2 = (add_ln703_729_reg_4897 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_836_fu_2655_p2 = (add_ln703_730_fu_2424_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_837_fu_2660_p2 = (add_ln703_732_reg_4902 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_838_fu_2664_p2 = (add_ln703_733_fu_2434_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_fu_248_p2 = (trunc_ln203_reg_3431 - tmp_2_reg_3437);

assign tmp_2_fu_92_p4 = {{data_V_read_int_reg[31:16]}};

assign trunc_ln203_fu_88_p1 = data_V_read_int_reg[15:0];

endmodule //dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;

reg   [15:0] data_31_V_read32_reg_4221;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter1_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter2_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter3_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter4_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter5_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter6_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter7_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter8_reg;
reg   [15:0] data_30_V_read31_reg_4250;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter1_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter2_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter3_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter4_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter5_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter6_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter7_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter8_reg;
reg   [15:0] data_29_V_read_7_reg_4279;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter1_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter2_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter3_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter4_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter5_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter6_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter7_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter8_reg;
reg   [15:0] data_28_V_read_7_reg_4313;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter1_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter2_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter3_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter4_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter5_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter6_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter7_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter8_reg;
reg   [15:0] data_27_V_read_8_reg_4342;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter1_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter2_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter3_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter4_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter5_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter6_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter7_reg;
reg   [15:0] data_26_V_read27_reg_4365;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter1_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter2_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter3_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter4_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter5_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter6_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter7_reg;
reg   [15:0] data_25_V_read26_reg_4391;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter1_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter2_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter3_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter4_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter5_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter6_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter7_reg;
reg   [15:0] data_24_V_read25_reg_4421;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter1_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter2_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter3_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter4_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter5_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter6_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter7_reg;
reg   [15:0] data_23_V_read24_reg_4451;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter1_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter2_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter3_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter4_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter5_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter6_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter7_reg;
reg   [15:0] data_22_V_read23_reg_4483;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter1_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter2_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter3_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter5_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter6_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter7_reg;
reg   [15:0] data_21_V_read22_reg_4512;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter1_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter2_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter3_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter4_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter5_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter6_reg;
reg   [15:0] data_20_V_read21_reg_4539;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter1_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter2_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter3_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter4_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter5_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter6_reg;
reg   [15:0] data_19_V_read_7_reg_4567;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter1_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter2_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter3_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter4_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter5_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter6_reg;
reg   [15:0] data_18_V_read_7_reg_4594;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter1_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter2_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter3_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter4_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter5_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter6_reg;
reg   [15:0] data_17_V_read_8_reg_4621;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter1_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter2_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter3_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter4_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter5_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter6_reg;
reg   [15:0] data_16_V_read17_reg_4650;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter1_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter2_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter3_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter4_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter5_reg;
reg   [15:0] data_15_V_read16_reg_4682;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter1_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter2_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter3_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter4_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter5_reg;
reg   [15:0] data_14_V_read15_reg_4714;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter1_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter2_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter3_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter4_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter5_reg;
reg   [15:0] data_13_V_read14_reg_4745;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter1_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter2_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter3_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter4_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter5_reg;
reg   [15:0] data_12_V_read13_reg_4778;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter1_reg;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter2_reg;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter3_reg;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter4_reg;
reg   [15:0] data_11_V_read12_reg_4808;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter1_reg;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter2_reg;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter3_reg;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter4_reg;
reg   [15:0] data_10_V_read11_reg_4832;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter1_reg;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter2_reg;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter3_reg;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter4_reg;
reg   [15:0] data_9_V_read_7_reg_4859;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter1_reg;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter2_reg;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter3_reg;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter4_reg;
reg   [15:0] data_8_V_read_7_reg_4887;
reg   [15:0] data_8_V_read_7_reg_4887_pp0_iter1_reg;
reg   [15:0] data_8_V_read_7_reg_4887_pp0_iter2_reg;
reg   [15:0] data_8_V_read_7_reg_4887_pp0_iter3_reg;
reg   [15:0] data_7_V_read_8_reg_4916;
reg   [15:0] data_7_V_read_8_reg_4916_pp0_iter1_reg;
reg   [15:0] data_7_V_read_8_reg_4916_pp0_iter2_reg;
reg   [15:0] data_7_V_read_8_reg_4916_pp0_iter3_reg;
reg   [15:0] data_6_V_read_8_reg_4944;
reg   [15:0] data_6_V_read_8_reg_4944_pp0_iter1_reg;
reg   [15:0] data_6_V_read_8_reg_4944_pp0_iter2_reg;
reg   [15:0] data_6_V_read_8_reg_4944_pp0_iter3_reg;
reg   [15:0] data_5_V_read_8_reg_4969;
reg   [15:0] data_5_V_read_8_reg_4969_pp0_iter1_reg;
reg   [15:0] data_5_V_read_8_reg_4969_pp0_iter2_reg;
reg   [15:0] data_5_V_read_8_reg_4969_pp0_iter3_reg;
reg   [15:0] data_4_V_read_9_reg_4998;
reg   [15:0] data_4_V_read_9_reg_4998_pp0_iter1_reg;
reg   [15:0] data_4_V_read_9_reg_4998_pp0_iter2_reg;
reg   [15:0] data_3_V_read_9_reg_5019;
reg   [15:0] data_3_V_read_9_reg_5019_pp0_iter1_reg;
reg   [15:0] data_3_V_read_9_reg_5019_pp0_iter2_reg;
reg   [15:0] data_2_V_read_9_reg_5035;
wire   [15:0] sub_ln703_fu_274_p2;
reg   [15:0] sub_ln703_reg_5046;
wire   [15:0] add_ln703_fu_280_p2;
reg   [15:0] add_ln703_reg_5052;
wire   [15:0] sub_ln703_73_fu_286_p2;
reg   [15:0] sub_ln703_73_reg_5059;
wire   [15:0] sub_ln703_74_fu_292_p2;
reg   [15:0] sub_ln703_74_reg_5065;
reg   [15:0] sub_ln703_74_reg_5065_pp0_iter2_reg;
wire   [15:0] sub_ln703_76_fu_300_p2;
reg   [15:0] sub_ln703_76_reg_5071;
reg   [15:0] sub_ln703_76_reg_5071_pp0_iter2_reg;
wire   [15:0] add_ln703_200_fu_304_p2;
reg   [15:0] add_ln703_200_reg_5077;
reg   [15:0] add_ln703_200_reg_5077_pp0_iter2_reg;
wire   [15:0] sub_ln703_77_fu_308_p2;
reg   [15:0] sub_ln703_77_reg_5084;
wire   [15:0] add_ln703_201_fu_312_p2;
reg   [15:0] add_ln703_201_reg_5090;
reg   [15:0] add_ln703_201_reg_5090_pp0_iter2_reg;
wire   [15:0] add_ln703_202_fu_316_p2;
reg   [15:0] add_ln703_202_reg_5096;
reg   [15:0] add_ln703_202_reg_5096_pp0_iter2_reg;
wire   [15:0] add_ln703_204_fu_320_p2;
reg   [15:0] add_ln703_204_reg_5101;
reg   [15:0] add_ln703_204_reg_5101_pp0_iter2_reg;
wire   [15:0] add_ln703_207_fu_325_p2;
reg   [15:0] add_ln703_207_reg_5107;
reg   [15:0] add_ln703_207_reg_5107_pp0_iter2_reg;
wire   [15:0] add_ln703_203_fu_329_p2;
reg   [15:0] add_ln703_203_reg_5113;
wire   [15:0] add_ln703_205_fu_333_p2;
reg   [15:0] add_ln703_205_reg_5119;
wire   [15:0] sub_ln703_79_fu_337_p2;
reg   [15:0] sub_ln703_79_reg_5125;
wire   [15:0] add_ln703_206_fu_341_p2;
reg   [15:0] add_ln703_206_reg_5131;
wire   [15:0] add_ln703_208_fu_345_p2;
reg   [15:0] add_ln703_208_reg_5137;
wire   [15:0] add_ln703_210_fu_349_p2;
reg   [15:0] add_ln703_210_reg_5143;
reg   [15:0] add_ln703_210_reg_5143_pp0_iter3_reg;
wire   [15:0] add_ln703_233_fu_353_p2;
reg   [15:0] add_ln703_233_reg_5149;
reg   [15:0] add_ln703_233_reg_5149_pp0_iter3_reg;
wire   [15:0] add_ln703_247_fu_357_p2;
reg   [15:0] add_ln703_247_reg_5159;
reg   [15:0] add_ln703_247_reg_5159_pp0_iter3_reg;
wire   [15:0] sub_ln703_89_fu_402_p2;
reg   [15:0] sub_ln703_89_reg_5166;
wire   [15:0] sub_ln703_91_fu_411_p2;
reg   [15:0] sub_ln703_91_reg_5172;
wire   [15:0] add_ln703_209_fu_416_p2;
reg   [15:0] add_ln703_209_reg_5178;
wire   [15:0] add_ln703_211_fu_420_p2;
reg   [15:0] add_ln703_211_reg_5184;
wire   [15:0] add_ln703_213_fu_429_p2;
reg   [15:0] add_ln703_213_reg_5189;
wire   [15:0] add_ln703_214_fu_433_p2;
reg   [15:0] add_ln703_214_reg_5194;
wire   [15:0] sub_ln703_93_fu_442_p2;
reg   [15:0] sub_ln703_93_reg_5200;
wire   [15:0] sub_ln703_94_fu_446_p2;
reg   [15:0] sub_ln703_94_reg_5205;
wire   [15:0] sub_ln703_96_fu_456_p2;
reg   [15:0] sub_ln703_96_reg_5210;
wire   [15:0] add_ln703_216_fu_461_p2;
reg   [15:0] add_ln703_216_reg_5215;
wire   [15:0] add_ln703_220_fu_484_p2;
reg   [15:0] add_ln703_220_reg_5221;
wire   [15:0] sub_ln703_105_fu_489_p2;
reg   [15:0] sub_ln703_105_reg_5226;
wire   [15:0] add_ln703_223_fu_507_p2;
reg   [15:0] add_ln703_223_reg_5231;
wire   [15:0] add_ln703_225_fu_513_p2;
reg   [15:0] add_ln703_225_reg_5237;
wire   [15:0] add_ln703_227_fu_522_p2;
reg   [15:0] add_ln703_227_reg_5242;
wire   [15:0] sub_ln703_113_fu_533_p2;
reg   [15:0] sub_ln703_113_reg_5247;
wire   [15:0] sub_ln703_114_fu_549_p2;
reg   [15:0] sub_ln703_114_reg_5253;
wire   [15:0] sub_ln703_117_fu_554_p2;
reg   [15:0] sub_ln703_117_reg_5259;
wire   [15:0] add_ln703_234_fu_564_p2;
reg   [15:0] add_ln703_234_reg_5264;
wire   [15:0] add_ln703_238_fu_569_p2;
reg   [15:0] add_ln703_238_reg_5269;
wire   [15:0] sub_ln703_126_fu_574_p2;
reg   [15:0] sub_ln703_126_reg_5274;
wire   [15:0] sub_ln703_129_fu_579_p2;
reg   [15:0] sub_ln703_129_reg_5279;
wire   [15:0] sub_ln703_133_fu_584_p2;
reg   [15:0] sub_ln703_133_reg_5284;
wire   [15:0] add_ln703_251_fu_589_p2;
reg   [15:0] add_ln703_251_reg_5289;
wire   [15:0] add_ln703_258_fu_593_p2;
reg   [15:0] add_ln703_258_reg_5295;
wire   [15:0] add_ln703_272_fu_597_p2;
reg   [15:0] add_ln703_272_reg_5304;
reg   [15:0] add_ln703_272_reg_5304_pp0_iter4_reg;
wire   [15:0] add_ln703_304_fu_601_p2;
reg   [15:0] add_ln703_304_reg_5314;
wire   [15:0] add_ln703_246_fu_787_p2;
reg   [15:0] add_ln703_246_reg_5320;
wire   [15:0] sub_ln703_138_fu_816_p2;
reg   [15:0] sub_ln703_138_reg_5325;
wire   [15:0] sub_ln703_141_fu_835_p2;
reg   [15:0] sub_ln703_141_reg_5330;
wire   [15:0] sub_ln703_143_fu_844_p2;
reg   [15:0] sub_ln703_143_reg_5335;
wire   [15:0] sub_ln703_144_fu_858_p2;
reg   [15:0] sub_ln703_144_reg_5340;
wire   [15:0] sub_ln703_145_fu_863_p2;
reg   [15:0] sub_ln703_145_reg_5345;
wire   [15:0] sub_ln703_149_fu_901_p2;
reg   [15:0] sub_ln703_149_reg_5350;
wire   [15:0] sub_ln703_154_fu_920_p2;
reg   [15:0] sub_ln703_154_reg_5355;
wire   [15:0] add_ln703_261_fu_955_p2;
reg   [15:0] add_ln703_261_reg_5360;
wire   [15:0] sub_ln703_161_fu_960_p2;
reg   [15:0] sub_ln703_161_reg_5365;
wire   [15:0] sub_ln703_162_fu_980_p2;
reg   [15:0] sub_ln703_162_reg_5370;
wire   [15:0] sub_ln703_166_fu_1000_p2;
reg   [15:0] sub_ln703_166_reg_5375;
wire   [15:0] sub_ln703_171_fu_1015_p2;
reg   [15:0] sub_ln703_171_reg_5380;
wire   [15:0] sub_ln703_173_fu_1025_p2;
reg   [15:0] sub_ln703_173_reg_5385;
wire   [15:0] sub_ln703_176_fu_1040_p2;
reg   [15:0] sub_ln703_176_reg_5390;
wire   [15:0] sub_ln703_180_fu_1045_p2;
reg   [15:0] sub_ln703_180_reg_5395;
wire   [15:0] sub_ln703_181_fu_1050_p2;
reg   [15:0] sub_ln703_181_reg_5400;
wire   [15:0] add_ln703_267_fu_1055_p2;
reg   [15:0] add_ln703_267_reg_5405;
wire   [15:0] sub_ln703_182_fu_1060_p2;
reg   [15:0] sub_ln703_182_reg_5410;
wire   [15:0] add_ln703_268_fu_1065_p2;
reg   [15:0] add_ln703_268_reg_5415;
wire   [15:0] add_ln703_274_fu_1089_p2;
reg   [15:0] add_ln703_274_reg_5420;
wire   [15:0] sub_ln703_185_fu_1095_p2;
reg   [15:0] sub_ln703_185_reg_5425;
wire   [15:0] add_ln703_276_fu_1100_p2;
reg   [15:0] add_ln703_276_reg_5430;
wire   [15:0] add_ln703_278_fu_1105_p2;
reg   [15:0] add_ln703_278_reg_5435;
wire   [15:0] sub_ln703_187_fu_1110_p2;
reg   [15:0] sub_ln703_187_reg_5440;
wire   [15:0] sub_ln703_189_fu_1115_p2;
reg   [15:0] sub_ln703_189_reg_5445;
wire   [15:0] sub_ln703_191_fu_1120_p2;
reg   [15:0] sub_ln703_191_reg_5450;
wire   [15:0] add_ln703_281_fu_1129_p2;
reg   [15:0] add_ln703_281_reg_5455;
wire   [15:0] add_ln703_283_fu_1140_p2;
reg   [15:0] add_ln703_283_reg_5460;
wire   [15:0] sub_ln703_198_fu_1146_p2;
reg   [15:0] sub_ln703_198_reg_5465;
wire   [15:0] sub_ln703_199_fu_1151_p2;
reg   [15:0] sub_ln703_199_reg_5470;
wire   [15:0] add_ln703_288_fu_1156_p2;
reg   [15:0] add_ln703_288_reg_5475;
wire   [15:0] add_ln703_309_fu_1179_p2;
reg   [15:0] add_ln703_309_reg_5484;
wire   [15:0] add_ln703_314_fu_1183_p2;
reg   [15:0] add_ln703_314_reg_5490;
wire   [15:0] add_ln703_316_fu_1187_p2;
reg   [15:0] add_ln703_316_reg_5496;
wire   [15:0] sub_ln703_246_fu_1193_p2;
reg   [15:0] sub_ln703_246_reg_5501;
wire   [15:0] add_ln703_323_fu_1198_p2;
reg   [15:0] add_ln703_323_reg_5506;
wire   [15:0] sub_ln703_200_fu_1326_p2;
reg   [15:0] sub_ln703_200_reg_5515;
wire   [15:0] sub_ln703_203_fu_1339_p2;
reg   [15:0] sub_ln703_203_reg_5520;
wire   [15:0] add_ln703_287_fu_1354_p2;
reg   [15:0] add_ln703_287_reg_5525;
wire   [15:0] add_ln703_291_fu_1371_p2;
reg   [15:0] add_ln703_291_reg_5530;
wire   [15:0] sub_ln703_207_fu_1384_p2;
reg   [15:0] sub_ln703_207_reg_5535;
wire   [15:0] sub_ln703_212_fu_1412_p2;
reg   [15:0] sub_ln703_212_reg_5540;
wire   [15:0] sub_ln703_215_fu_1441_p2;
reg   [15:0] sub_ln703_215_reg_5545;
wire   [15:0] add_ln703_301_fu_1494_p2;
reg   [15:0] add_ln703_301_reg_5550;
wire   [15:0] add_ln703_307_fu_1504_p2;
reg   [15:0] add_ln703_307_reg_5555;
wire   [15:0] sub_ln703_229_fu_1518_p2;
reg   [15:0] sub_ln703_229_reg_5560;
wire   [15:0] sub_ln703_237_fu_1571_p2;
reg   [15:0] sub_ln703_237_reg_5565;
wire   [15:0] sub_ln703_238_fu_1576_p2;
reg   [15:0] sub_ln703_238_reg_5570;
wire   [15:0] sub_ln703_252_fu_1616_p2;
reg   [15:0] sub_ln703_252_reg_5575;
wire   [15:0] sub_ln703_253_fu_1621_p2;
reg   [15:0] sub_ln703_253_reg_5580;
wire   [15:0] sub_ln703_254_fu_1626_p2;
reg   [15:0] sub_ln703_254_reg_5585;
wire   [15:0] add_ln703_321_fu_1636_p2;
reg   [15:0] add_ln703_321_reg_5590;
wire   [15:0] sub_ln703_257_fu_1641_p2;
reg   [15:0] sub_ln703_257_reg_5595;
wire   [15:0] sub_ln703_261_fu_1646_p2;
reg   [15:0] sub_ln703_261_reg_5600;
wire   [15:0] sub_ln703_262_fu_1651_p2;
reg   [15:0] sub_ln703_262_reg_5605;
wire   [15:0] sub_ln703_263_fu_1671_p2;
reg   [15:0] sub_ln703_263_reg_5610;
wire   [15:0] sub_ln703_265_fu_1676_p2;
reg   [15:0] sub_ln703_265_reg_5615;
wire   [15:0] sub_ln703_266_fu_1681_p2;
reg   [15:0] sub_ln703_266_reg_5620;
wire   [15:0] add_ln703_326_fu_1686_p2;
reg   [15:0] add_ln703_326_reg_5625;
wire   [15:0] sub_ln703_270_fu_1695_p2;
reg   [15:0] sub_ln703_270_reg_5630;
wire   [15:0] sub_ln703_272_fu_1700_p2;
reg   [15:0] sub_ln703_272_reg_5635;
wire   [15:0] add_ln703_330_fu_1710_p2;
reg   [15:0] add_ln703_330_reg_5640;
wire   [15:0] add_ln703_335_fu_1730_p2;
reg   [15:0] add_ln703_335_reg_5645;
wire   [15:0] sub_ln703_278_fu_1735_p2;
reg   [15:0] sub_ln703_278_reg_5650;
wire   [15:0] add_ln703_339_fu_1740_p2;
reg   [15:0] add_ln703_339_reg_5655;
wire   [15:0] add_ln703_343_fu_1745_p2;
reg   [15:0] add_ln703_343_reg_5660;
wire   [15:0] sub_ln703_289_fu_1750_p2;
reg   [15:0] sub_ln703_289_reg_5665;
wire   [15:0] sub_ln703_290_fu_1755_p2;
reg   [15:0] sub_ln703_290_reg_5670;
wire   [15:0] add_ln703_347_fu_1760_p2;
reg   [15:0] add_ln703_347_reg_5675;
wire   [15:0] add_ln703_357_fu_1764_p2;
reg   [15:0] add_ln703_357_reg_5683;
reg   [15:0] add_ln703_357_reg_5683_pp0_iter6_reg;
wire   [15:0] add_ln703_371_fu_1768_p2;
reg   [15:0] add_ln703_371_reg_5691;
wire   [15:0] add_ln703_384_fu_1772_p2;
reg   [15:0] add_ln703_384_reg_5701;
reg   [15:0] add_ln703_384_reg_5701_pp0_iter6_reg;
wire   [15:0] add_ln703_394_fu_1776_p2;
reg   [15:0] add_ln703_394_reg_5710;
reg   [15:0] add_ln703_394_reg_5710_pp0_iter6_reg;
wire   [15:0] add_ln703_404_fu_1780_p2;
reg   [15:0] add_ln703_404_reg_5718;
reg   [15:0] add_ln703_404_reg_5718_pp0_iter6_reg;
wire   [15:0] sub_ln703_276_fu_1918_p2;
reg   [15:0] sub_ln703_276_reg_5728;
wire   [15:0] sub_ln703_283_fu_1975_p2;
reg   [15:0] sub_ln703_283_reg_5733;
wire   [15:0] sub_ln703_288_fu_2003_p2;
reg   [15:0] sub_ln703_288_reg_5738;
wire   [15:0] add_ln703_353_fu_2060_p2;
reg   [15:0] add_ln703_353_reg_5743;
wire   [15:0] sub_ln703_300_fu_2075_p2;
reg   [15:0] sub_ln703_300_reg_5748;
wire   [15:0] add_ln703_354_fu_2080_p2;
reg   [15:0] add_ln703_354_reg_5753;
wire   [15:0] sub_ln703_302_fu_2089_p2;
reg   [15:0] sub_ln703_302_reg_5758;
wire   [15:0] sub_ln703_304_fu_2099_p2;
reg   [15:0] sub_ln703_304_reg_5763;
wire   [15:0] add_ln703_359_fu_2127_p2;
reg   [15:0] add_ln703_359_reg_5768;
wire   [15:0] sub_ln703_309_fu_2148_p2;
reg   [15:0] sub_ln703_309_reg_5773;
wire   [15:0] sub_ln703_311_fu_2173_p2;
reg   [15:0] sub_ln703_311_reg_5778;
wire   [15:0] sub_ln703_318_fu_2203_p2;
reg   [15:0] sub_ln703_318_reg_5783;
wire   [15:0] sub_ln703_321_fu_2218_p2;
reg   [15:0] sub_ln703_321_reg_5788;
wire   [15:0] add_ln703_372_fu_2228_p2;
reg   [15:0] add_ln703_372_reg_5793;
wire   [15:0] sub_ln703_323_fu_2233_p2;
reg   [15:0] sub_ln703_323_reg_5798;
wire   [15:0] sub_ln703_324_fu_2238_p2;
reg   [15:0] sub_ln703_324_reg_5803;
wire   [15:0] sub_ln703_325_fu_2243_p2;
reg   [15:0] sub_ln703_325_reg_5808;
wire   [15:0] sub_ln703_327_fu_2248_p2;
reg   [15:0] sub_ln703_327_reg_5813;
wire   [15:0] sub_ln703_328_fu_2253_p2;
reg   [15:0] sub_ln703_328_reg_5818;
wire   [15:0] sub_ln703_331_fu_2258_p2;
reg   [15:0] sub_ln703_331_reg_5823;
wire   [15:0] sub_ln703_332_fu_2273_p2;
reg   [15:0] sub_ln703_332_reg_5828;
wire   [15:0] add_ln703_377_fu_2283_p2;
reg   [15:0] add_ln703_377_reg_5833;
wire   [15:0] add_ln703_379_fu_2292_p2;
reg   [15:0] add_ln703_379_reg_5838;
wire   [15:0] sub_ln703_335_fu_2302_p2;
reg   [15:0] sub_ln703_335_reg_5843;
wire   [15:0] add_ln703_381_fu_2307_p2;
reg   [15:0] add_ln703_381_reg_5848;
wire   [15:0] sub_ln703_343_fu_2312_p2;
reg   [15:0] sub_ln703_343_reg_5853;
wire   [15:0] add_ln703_390_fu_2326_p2;
reg   [15:0] add_ln703_390_reg_5858;
wire   [15:0] sub_ln703_346_fu_2332_p2;
reg   [15:0] sub_ln703_346_reg_5863;
wire   [15:0] add_ln703_400_fu_2346_p2;
reg   [15:0] add_ln703_400_reg_5868;
wire   [15:0] add_ln703_413_fu_2361_p2;
reg   [15:0] add_ln703_413_reg_5873;
wire   [15:0] add_ln703_415_fu_2372_p2;
reg   [15:0] add_ln703_415_reg_5878;
wire   [15:0] add_ln703_427_fu_2383_p2;
reg   [15:0] add_ln703_427_reg_5883;
wire   [15:0] add_ln703_428_fu_2389_p2;
reg   [15:0] add_ln703_428_reg_5888;
wire   [15:0] add_ln703_435_fu_2393_p2;
reg   [15:0] add_ln703_435_reg_5894;
wire   [15:0] add_ln703_446_fu_2397_p2;
reg   [15:0] add_ln703_446_reg_5901;
wire   [15:0] add_ln703_462_fu_2401_p2;
reg   [15:0] add_ln703_462_reg_5909;
reg   [15:0] add_ln703_462_reg_5909_pp0_iter7_reg;
reg   [15:0] add_ln703_462_reg_5909_pp0_iter8_reg;
wire   [15:0] sub_ln703_356_fu_2603_p2;
reg   [15:0] sub_ln703_356_reg_5921;
wire   [15:0] sub_ln703_357_fu_2608_p2;
reg   [15:0] sub_ln703_357_reg_5926;
wire   [15:0] add_ln703_402_fu_2631_p2;
reg   [15:0] add_ln703_402_reg_5931;
wire   [15:0] sub_ln703_361_fu_2636_p2;
reg   [15:0] sub_ln703_361_reg_5936;
wire   [15:0] sub_ln703_366_fu_2684_p2;
reg   [15:0] sub_ln703_366_reg_5941;
wire   [15:0] sub_ln703_369_fu_2699_p2;
reg   [15:0] sub_ln703_369_reg_5946;
wire   [15:0] add_ln703_410_fu_2709_p2;
reg   [15:0] add_ln703_410_reg_5951;
wire   [15:0] sub_ln703_374_fu_2728_p2;
reg   [15:0] sub_ln703_374_reg_5956;
wire   [15:0] add_ln703_418_fu_2741_p2;
reg   [15:0] add_ln703_418_reg_5961;
wire   [15:0] sub_ln703_375_fu_2747_p2;
reg   [15:0] sub_ln703_375_reg_5966;
wire   [15:0] sub_ln703_379_fu_2781_p2;
reg   [15:0] sub_ln703_379_reg_5971;
wire   [15:0] sub_ln703_381_fu_2791_p2;
reg   [15:0] sub_ln703_381_reg_5976;
wire   [15:0] add_ln703_424_fu_2806_p2;
reg   [15:0] add_ln703_424_reg_5981;
wire   [15:0] sub_ln703_385_fu_2811_p2;
reg   [15:0] sub_ln703_385_reg_5986;
wire   [15:0] sub_ln703_386_fu_2816_p2;
reg   [15:0] sub_ln703_386_reg_5991;
wire   [15:0] sub_ln703_389_fu_2839_p2;
reg   [15:0] sub_ln703_389_reg_5996;
wire   [15:0] sub_ln703_392_fu_2848_p2;
reg   [15:0] sub_ln703_392_reg_6001;
wire   [15:0] sub_ln703_397_fu_2863_p2;
reg   [15:0] sub_ln703_397_reg_6006;
wire   [15:0] add_ln703_434_fu_2873_p2;
reg   [15:0] add_ln703_434_reg_6011;
wire   [15:0] sub_ln703_402_fu_2878_p2;
reg   [15:0] sub_ln703_402_reg_6016;
wire   [15:0] add_ln703_436_fu_2883_p2;
reg   [15:0] add_ln703_436_reg_6021;
wire   [15:0] sub_ln703_408_fu_2893_p2;
reg   [15:0] sub_ln703_408_reg_6026;
wire   [15:0] sub_ln703_409_fu_2898_p2;
reg   [15:0] sub_ln703_409_reg_6031;
wire   [15:0] sub_ln703_411_fu_2903_p2;
reg   [15:0] sub_ln703_411_reg_6036;
wire   [15:0] add_ln703_442_fu_2917_p2;
reg   [15:0] add_ln703_442_reg_6041;
wire   [15:0] sub_ln703_416_fu_2923_p2;
reg   [15:0] sub_ln703_416_reg_6046;
wire   [15:0] add_ln703_444_fu_2928_p2;
reg   [15:0] add_ln703_444_reg_6051;
wire   [15:0] add_ln703_447_fu_2933_p2;
reg   [15:0] add_ln703_447_reg_6056;
wire   [15:0] sub_ln703_426_fu_2938_p2;
reg   [15:0] sub_ln703_426_reg_6061;
wire   [15:0] add_ln703_451_fu_2943_p2;
reg   [15:0] add_ln703_451_reg_6066;
reg   [15:0] add_ln703_451_reg_6066_pp0_iter8_reg;
wire   [15:0] add_ln703_480_fu_2961_p2;
reg   [15:0] add_ln703_480_reg_6072;
reg   [15:0] add_ln703_480_reg_6072_pp0_iter8_reg;
wire   [15:0] add_ln703_482_fu_2967_p2;
reg   [15:0] add_ln703_482_reg_6077;
wire   [15:0] add_ln703_491_fu_2971_p2;
reg   [15:0] add_ln703_491_reg_6087;
reg   [15:0] add_ln703_491_reg_6087_pp0_iter8_reg;
wire   [15:0] add_ln703_509_fu_2976_p2;
reg   [15:0] add_ln703_509_reg_6092;
reg   [15:0] add_ln703_509_reg_6092_pp0_iter8_reg;
wire   [15:0] add_ln703_516_fu_2980_p2;
reg   [15:0] add_ln703_516_reg_6103;
reg   [15:0] add_ln703_516_reg_6103_pp0_iter8_reg;
wire   [15:0] sub_ln703_428_fu_3163_p2;
reg   [15:0] sub_ln703_428_reg_6108;
wire   [15:0] sub_ln703_434_fu_3199_p2;
reg   [15:0] sub_ln703_434_reg_6113;
wire   [15:0] sub_ln703_448_fu_3308_p2;
reg   [15:0] sub_ln703_448_reg_6118;
wire   [15:0] sub_ln703_450_fu_3318_p2;
reg   [15:0] sub_ln703_450_reg_6123;
wire   [15:0] add_ln703_463_fu_3328_p2;
reg   [15:0] add_ln703_463_reg_6128;
wire   [15:0] add_ln703_464_fu_3333_p2;
reg   [15:0] add_ln703_464_reg_6133;
wire   [15:0] add_ln703_465_fu_3338_p2;
reg   [15:0] add_ln703_465_reg_6138;
wire   [15:0] sub_ln703_451_fu_3343_p2;
reg   [15:0] sub_ln703_451_reg_6143;
wire   [15:0] sub_ln703_452_fu_3348_p2;
reg   [15:0] sub_ln703_452_reg_6148;
wire   [15:0] sub_ln703_453_fu_3353_p2;
reg   [15:0] sub_ln703_453_reg_6153;
wire   [15:0] add_ln703_467_fu_3363_p2;
reg   [15:0] add_ln703_467_reg_6158;
wire   [15:0] sub_ln703_454_fu_3368_p2;
reg   [15:0] sub_ln703_454_reg_6163;
wire   [15:0] sub_ln703_455_fu_3373_p2;
reg   [15:0] sub_ln703_455_reg_6168;
wire   [15:0] add_ln703_468_fu_3378_p2;
reg   [15:0] add_ln703_468_reg_6173;
wire   [15:0] sub_ln703_456_fu_3388_p2;
reg   [15:0] sub_ln703_456_reg_6178;
wire   [15:0] sub_ln703_457_fu_3393_p2;
reg   [15:0] sub_ln703_457_reg_6183;
wire   [15:0] add_ln703_471_fu_3403_p2;
reg   [15:0] add_ln703_471_reg_6188;
wire   [15:0] sub_ln703_458_fu_3408_p2;
reg   [15:0] sub_ln703_458_reg_6193;
wire   [15:0] sub_ln703_459_fu_3418_p2;
reg   [15:0] sub_ln703_459_reg_6198;
wire   [15:0] add_ln703_475_fu_3432_p2;
reg   [15:0] add_ln703_475_reg_6203;
wire   [15:0] sub_ln703_461_fu_3438_p2;
reg   [15:0] sub_ln703_461_reg_6208;
wire   [15:0] add_ln703_483_fu_3448_p2;
reg   [15:0] add_ln703_483_reg_6213;
wire   [15:0] sub_ln703_469_fu_3463_p2;
reg   [15:0] sub_ln703_469_reg_6218;
wire   [15:0] add_ln703_492_fu_3478_p2;
reg   [15:0] add_ln703_492_reg_6223;
wire   [15:0] sub_ln703_474_fu_3482_p2;
reg   [15:0] sub_ln703_474_reg_6229;
wire   [15:0] add_ln703_496_fu_3497_p2;
reg   [15:0] add_ln703_496_reg_6234;
wire   [15:0] add_ln703_497_fu_3501_p2;
reg   [15:0] add_ln703_497_reg_6239;
wire   [15:0] sub_ln703_486_fu_3507_p2;
reg   [15:0] sub_ln703_486_reg_6244;
wire   [15:0] sub_ln703_487_fu_3512_p2;
reg   [15:0] sub_ln703_487_reg_6249;
wire   [15:0] sub_ln703_491_fu_3517_p2;
reg   [15:0] sub_ln703_491_reg_6254;
wire   [15:0] sub_ln703_500_fu_3522_p2;
reg   [15:0] sub_ln703_500_reg_6259;
wire   [15:0] add_ln703_510_fu_3527_p2;
reg   [15:0] add_ln703_510_reg_6264;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_75_fu_296_p2;
wire   [15:0] sub_ln703_78_fu_361_p2;
wire   [15:0] sub_ln703_80_fu_365_p2;
wire   [15:0] sub_ln703_81_fu_369_p2;
wire   [15:0] sub_ln703_82_fu_373_p2;
wire   [15:0] sub_ln703_84_fu_381_p2;
wire   [15:0] sub_ln703_86_fu_389_p2;
wire   [15:0] sub_ln703_87_fu_393_p2;
wire   [15:0] sub_ln703_88_fu_398_p2;
wire   [15:0] sub_ln703_90_fu_406_p2;
wire   [15:0] add_ln703_212_fu_425_p2;
wire   [15:0] sub_ln703_92_fu_437_p2;
wire   [15:0] add_ln703_222_fu_503_p2;
wire   [15:0] sub_ln703_85_fu_385_p2;
wire   [15:0] sub_ln703_98_fu_466_p2;
wire   [15:0] add_ln703_226_fu_518_p2;
wire   [15:0] add_ln703_217_fu_470_p2;
wire   [15:0] add_ln703_218_fu_474_p2;
wire   [15:0] sub_ln703_83_fu_377_p2;
wire   [15:0] add_ln703_230_fu_538_p2;
wire   [15:0] add_ln703_219_fu_479_p2;
wire   [15:0] sub_ln703_106_fu_494_p2;
wire   [15:0] add_ln703_221_fu_499_p2;
wire   [15:0] sub_ln703_95_fu_451_p2;
wire   [15:0] sub_ln703_112_fu_528_p2;
wire   [15:0] add_ln703_231_fu_543_p2;
wire   [15:0] sub_ln703_118_fu_559_p2;
wire   [15:0] add_ln703_215_fu_605_p2;
wire   [15:0] sub_ln703_97_fu_609_p2;
wire   [15:0] sub_ln703_99_fu_613_p2;
wire   [15:0] sub_ln703_100_fu_617_p2;
wire   [15:0] sub_ln703_101_fu_621_p2;
wire   [15:0] sub_ln703_103_fu_629_p2;
wire   [15:0] sub_ln703_108_fu_641_p2;
wire   [15:0] add_ln703_224_fu_645_p2;
wire   [15:0] sub_ln703_110_fu_654_p2;
wire   [15:0] sub_ln703_111_fu_658_p2;
wire   [15:0] add_ln703_228_fu_663_p2;
wire   [15:0] add_ln703_229_fu_668_p2;
wire   [15:0] add_ln703_232_fu_673_p2;
wire   [15:0] sub_ln703_102_fu_625_p2;
wire   [15:0] sub_ln703_115_fu_678_p2;
wire   [15:0] sub_ln703_116_fu_683_p2;
wire   [15:0] sub_ln703_107_fu_637_p2;
wire   [15:0] add_ln703_243_fu_774_p2;
wire   [15:0] sub_ln703_119_fu_687_p2;
wire   [15:0] sub_ln703_121_fu_696_p2;
wire   [15:0] sub_ln703_109_fu_649_p2;
wire   [15:0] add_ln703_235_fu_701_p2;
wire   [15:0] sub_ln703_122_fu_705_p2;
wire   [15:0] add_ln703_236_fu_710_p2;
wire   [15:0] add_ln703_237_fu_715_p2;
wire   [15:0] sub_ln703_123_fu_719_p2;
wire   [15:0] sub_ln703_125_fu_727_p2;
wire   [15:0] sub_ln703_128_fu_736_p2;
wire   [15:0] add_ln703_250_fu_849_p2;
wire   [15:0] add_ln703_239_fu_750_p2;
wire   [15:0] add_ln703_240_fu_755_p2;
wire   [15:0] sub_ln703_132_fu_760_p2;
wire   [15:0] add_ln703_253_fu_873_p2;
wire   [15:0] add_ln703_241_fu_765_p2;
wire   [15:0] add_ln703_255_fu_887_p2;
wire   [15:0] add_ln703_242_fu_769_p2;
wire   [15:0] add_ln703_244_fu_778_p2;
wire   [15:0] add_ln703_245_fu_783_p2;
wire   [15:0] sub_ln703_134_fu_792_p2;
wire   [15:0] add_ln703_248_fu_801_p2;
wire   [15:0] sub_ln703_139_fu_821_p2;
wire   [15:0] sub_ln703_140_fu_826_p2;
wire   [15:0] add_ln703_249_fu_830_p2;
wire   [15:0] sub_ln703_124_fu_723_p2;
wire   [15:0] sub_ln703_142_fu_840_p2;
wire   [15:0] sub_ln703_127_fu_732_p2;
wire   [15:0] sub_ln703_131_fu_745_p2;
wire   [15:0] add_ln703_252_fu_853_p2;
wire   [15:0] sub_ln703_104_fu_633_p2;
wire   [15:0] add_ln703_263_fu_970_p2;
wire   [15:0] add_ln703_262_fu_965_p2;
wire   [15:0] sub_ln703_146_fu_868_p2;
wire   [15:0] add_ln703_254_fu_877_p2;
wire   [15:0] sub_ln703_147_fu_882_p2;
wire   [15:0] add_ln703_256_fu_891_p2;
wire   [15:0] sub_ln703_148_fu_896_p2;
wire   [15:0] sub_ln703_151_fu_911_p2;
wire   [15:0] sub_ln703_153_fu_915_p2;
wire   [15:0] add_ln703_257_fu_925_p2;
wire   [15:0] sub_ln703_156_fu_930_p2;
wire   [15:0] sub_ln703_157_fu_935_p2;
wire   [15:0] add_ln703_259_fu_940_p2;
wire   [15:0] sub_ln703_159_fu_945_p2;
wire   [15:0] add_ln703_260_fu_950_p2;
wire   [15:0] add_ln703_264_fu_974_p2;
wire   [15:0] sub_ln703_163_fu_985_p2;
wire   [15:0] sub_ln703_164_fu_990_p2;
wire   [15:0] sub_ln703_165_fu_995_p2;
wire   [15:0] sub_ln703_150_fu_906_p2;
wire   [15:0] sub_ln703_168_fu_1005_p2;
wire   [15:0] sub_ln703_120_fu_691_p2;
wire   [15:0] add_ln703_273_fu_1085_p2;
wire   [15:0] add_ln703_271_fu_1080_p2;
wire   [15:0] add_ln703_265_fu_1010_p2;
wire   [15:0] sub_ln703_136_fu_806_p2;
wire   [15:0] sub_ln703_137_fu_811_p2;
wire   [15:0] sub_ln703_172_fu_1020_p2;
wire   [15:0] sub_ln703_174_fu_1030_p2;
wire   [15:0] sub_ln703_175_fu_1035_p2;
wire   [15:0] add_ln703_280_fu_1125_p2;
wire   [15:0] sub_ln703_130_fu_741_p2;
wire   [15:0] add_ln703_282_fu_1135_p2;
wire   [15:0] add_ln703_269_fu_1069_p2;
wire   [15:0] sub_ln703_184_fu_1075_p2;
wire   [15:0] add_ln703_302_fu_1160_p2;
wire   [15:0] add_ln703_305_fu_1169_p2;
wire   [15:0] add_ln703_303_fu_1164_p2;
wire   [15:0] sub_ln703_135_fu_796_p2;
wire   [15:0] add_ln703_306_fu_1173_p2;
wire   [15:0] sub_ln703_152_fu_1202_p2;
wire   [15:0] sub_ln703_155_fu_1206_p2;
wire   [15:0] sub_ln703_158_fu_1210_p2;
wire   [15:0] sub_ln703_160_fu_1214_p2;
wire   [15:0] sub_ln703_167_fu_1218_p2;
wire   [15:0] sub_ln703_169_fu_1222_p2;
wire   [15:0] sub_ln703_170_fu_1227_p2;
wire   [15:0] add_ln703_266_fu_1232_p2;
wire   [15:0] sub_ln703_177_fu_1237_p2;
wire   [15:0] sub_ln703_179_fu_1246_p2;
wire   [15:0] add_ln703_284_fu_1296_p2;
wire   [15:0] sub_ln703_183_fu_1250_p2;
wire   [15:0] add_ln703_270_fu_1255_p2;
wire   [15:0] add_ln703_275_fu_1260_p2;
wire   [15:0] add_ln703_277_fu_1264_p2;
wire   [15:0] add_ln703_279_fu_1268_p2;
wire   [15:0] sub_ln703_186_fu_1272_p2;
wire   [15:0] sub_ln703_190_fu_1281_p2;
wire   [15:0] sub_ln703_192_fu_1286_p2;
wire   [15:0] sub_ln703_178_fu_1242_p2;
wire   [15:0] sub_ln703_193_fu_1291_p2;
wire   [15:0] add_ln703_285_fu_1300_p2;
wire   [15:0] add_ln703_286_fu_1305_p2;
wire   [15:0] sub_ln703_194_fu_1309_p2;
wire   [15:0] sub_ln703_195_fu_1313_p2;
wire   [15:0] sub_ln703_196_fu_1317_p2;
wire   [15:0] add_ln703_296_fu_1432_p2;
wire   [15:0] sub_ln703_197_fu_1321_p2;
wire   [15:0] sub_ln703_202_fu_1335_p2;
wire   [15:0] sub_ln703_204_fu_1344_p2;
wire   [15:0] sub_ln703_205_fu_1349_p2;
wire   [15:0] add_ln703_289_fu_1359_p2;
wire   [15:0] sub_ln703_206_fu_1363_p2;
wire   [15:0] add_ln703_290_fu_1367_p2;
wire   [15:0] add_ln703_292_fu_1376_p2;
wire   [15:0] add_ln703_293_fu_1380_p2;
wire   [15:0] sub_ln703_208_fu_1389_p2;
wire   [15:0] add_ln703_294_fu_1397_p2;
wire   [15:0] sub_ln703_210_fu_1402_p2;
wire   [15:0] add_ln703_308_fu_1509_p2;
wire   [15:0] sub_ln703_211_fu_1407_p2;
wire   [15:0] add_ln703_311_fu_1523_p2;
wire   [15:0] sub_ln703_213_fu_1417_p2;
wire   [15:0] add_ln703_295_fu_1427_p2;
wire   [15:0] add_ln703_297_fu_1436_p2;
wire   [15:0] sub_ln703_217_fu_1450_p2;
wire   [15:0] sub_ln703_201_fu_1331_p2;
wire   [15:0] add_ln703_298_fu_1454_p2;
wire   [15:0] add_ln703_317_fu_1562_p2;
wire   [15:0] sub_ln703_220_fu_1459_p2;
wire   [15:0] add_ln703_299_fu_1464_p2;
wire   [15:0] sub_ln703_222_fu_1469_p2;
wire   [15:0] add_ln703_300_fu_1474_p2;
wire   [15:0] sub_ln703_223_fu_1479_p2;
wire   [15:0] sub_ln703_225_fu_1484_p2;
wire   [15:0] sub_ln703_226_fu_1489_p2;
wire   [15:0] add_ln703_310_fu_1513_p2;
wire   [15:0] add_ln703_312_fu_1527_p2;
wire   [15:0] add_ln703_313_fu_1532_p2;
wire   [15:0] sub_ln703_231_fu_1537_p2;
wire   [15:0] sub_ln703_232_fu_1542_p2;
wire   [15:0] add_ln703_315_fu_1552_p2;
wire   [15:0] sub_ln703_236_fu_1557_p2;
wire   [15:0] add_ln703_318_fu_1566_p2;
wire   [15:0] sub_ln703_240_fu_1581_p2;
wire   [15:0] sub_ln703_241_fu_1586_p2;
wire   [15:0] sub_ln703_188_fu_1277_p2;
wire   [15:0] add_ln703_324_fu_1661_p2;
wire   [15:0] add_ln703_322_fu_1656_p2;
wire   [15:0] add_ln703_319_fu_1591_p2;
wire   [15:0] sub_ln703_242_fu_1596_p2;
wire   [15:0] sub_ln703_243_fu_1601_p2;
wire   [15:0] sub_ln703_228_fu_1499_p2;
wire   [15:0] sub_ln703_248_fu_1606_p2;
wire   [15:0] sub_ln703_251_fu_1611_p2;
wire   [15:0] sub_ln703_214_fu_1422_p2;
wire   [15:0] add_ln703_329_fu_1705_p2;
wire   [15:0] sub_ln703_216_fu_1446_p2;
wire   [15:0] add_ln703_332_fu_1715_p2;
wire   [15:0] sub_ln703_234_fu_1547_p2;
wire   [15:0] sub_ln703_256_fu_1631_p2;
wire   [15:0] add_ln703_325_fu_1665_p2;
wire   [15:0] sub_ln703_209_fu_1393_p2;
wire   [15:0] sub_ln703_268_fu_1691_p2;
wire   [15:0] add_ln703_333_fu_1720_p2;
wire   [15:0] add_ln703_334_fu_1725_p2;
wire   [15:0] sub_ln703_218_fu_1784_p2;
wire   [15:0] sub_ln703_221_fu_1792_p2;
wire   [15:0] sub_ln703_224_fu_1796_p2;
wire   [15:0] sub_ln703_227_fu_1800_p2;
wire   [15:0] sub_ln703_230_fu_1804_p2;
wire   [15:0] sub_ln703_233_fu_1808_p2;
wire   [15:0] sub_ln703_239_fu_1817_p2;
wire   [15:0] add_ln703_320_fu_1822_p2;
wire   [15:0] sub_ln703_245_fu_1832_p2;
wire   [15:0] sub_ln703_247_fu_1836_p2;
wire   [15:0] sub_ln703_249_fu_1840_p2;
wire   [15:0] sub_ln703_250_fu_1844_p2;
wire   [15:0] sub_ln703_255_fu_1849_p2;
wire   [15:0] sub_ln703_258_fu_1854_p2;
wire   [15:0] sub_ln703_260_fu_1862_p2;
wire   [15:0] add_ln703_340_fu_1943_p2;
wire   [15:0] add_ln703_341_fu_1947_p2;
wire   [15:0] sub_ln703_269_fu_1877_p2;
wire   [15:0] sub_ln703_271_fu_1882_p2;
wire   [15:0] add_ln703_327_fu_1887_p2;
wire   [15:0] add_ln703_328_fu_1892_p2;
wire   [15:0] sub_ln703_273_fu_1896_p2;
wire   [15:0] add_ln703_331_fu_1900_p2;
wire   [15:0] sub_ln703_274_fu_1904_p2;
wire   [15:0] sub_ln703_275_fu_1909_p2;
wire   [15:0] sub_ln703_219_fu_1788_p2;
wire   [15:0] add_ln703_350_fu_2026_p2;
wire   [15:0] add_ln703_349_fu_2021_p2;
wire   [15:0] add_ln703_336_fu_1913_p2;
wire   [15:0] add_ln703_337_fu_1923_p2;
wire   [15:0] sub_ln703_277_fu_1927_p2;
wire   [15:0] sub_ln703_279_fu_1931_p2;
wire   [15:0] sub_ln703_264_fu_1867_p2;
wire   [15:0] sub_ln703_280_fu_1935_p2;
wire   [15:0] add_ln703_338_fu_1939_p2;
wire   [15:0] add_ln703_342_fu_1952_p2;
wire   [15:0] sub_ln703_281_fu_1957_p2;
wire   [15:0] sub_ln703_282_fu_1961_p2;
wire   [15:0] add_ln703_344_fu_1966_p2;
wire   [15:0] add_ln703_345_fu_1970_p2;
wire   [15:0] sub_ln703_286_fu_1989_p2;
wire   [15:0] add_ln703_346_fu_1993_p2;
wire   [15:0] sub_ln703_235_fu_1812_p2;
wire   [15:0] add_ln703_358_fu_2123_p2;
wire   [15:0] add_ln703_356_fu_2118_p2;
wire   [15:0] sub_ln703_291_fu_2008_p2;
wire   [15:0] sub_ln703_292_fu_2012_p2;
wire   [15:0] add_ln703_348_fu_2017_p2;
wire   [15:0] add_ln703_351_fu_2030_p2;
wire   [15:0] sub_ln703_259_fu_1858_p2;
wire   [15:0] add_ln703_361_fu_2153_p2;
wire   [15:0] sub_ln703_295_fu_2041_p2;
wire   [15:0] sub_ln703_296_fu_2046_p2;
wire   [15:0] add_ln703_352_fu_2051_p2;
wire   [15:0] sub_ln703_297_fu_2055_p2;
wire   [15:0] sub_ln703_298_fu_2065_p2;
wire   [15:0] sub_ln703_301_fu_2085_p2;
wire   [15:0] sub_ln703_303_fu_2094_p2;
wire   [15:0] sub_ln703_305_fu_2104_p2;
wire   [15:0] sub_ln703_306_fu_2109_p2;
wire   [15:0] add_ln703_355_fu_2114_p2;
wire   [15:0] sub_ln703_307_fu_2133_p2;
wire   [15:0] add_ln703_360_fu_2138_p2;
wire   [15:0] sub_ln703_308_fu_2143_p2;
wire   [15:0] sub_ln703_293_fu_2036_p2;
wire   [15:0] add_ln703_362_fu_2158_p2;
wire   [15:0] add_ln703_363_fu_2163_p2;
wire   [15:0] sub_ln703_310_fu_2168_p2;
wire   [15:0] add_ln703_364_fu_2178_p2;
wire   [15:0] add_ln703_365_fu_2183_p2;
wire   [15:0] add_ln703_366_fu_2193_p2;
wire   [15:0] sub_ln703_284_fu_1980_p2;
wire   [15:0] add_ln703_374_fu_2263_p2;
wire   [15:0] add_ln703_367_fu_2198_p2;
wire   [15:0] sub_ln703_287_fu_1998_p2;
wire   [15:0] add_ln703_376_fu_2278_p2;
wire   [15:0] add_ln703_378_fu_2288_p2;
wire   [15:0] sub_ln703_319_fu_2208_p2;
wire   [15:0] add_ln703_369_fu_2213_p2;
wire   [15:0] sub_ln703_322_fu_2223_p2;
wire   [15:0] add_ln703_375_fu_2268_p2;
wire   [15:0] sub_ln703_285_fu_1984_p2;
wire   [15:0] add_ln703_389_fu_2322_p2;
wire   [15:0] add_ln703_388_fu_2317_p2;
wire   [15:0] add_ln703_380_fu_2297_p2;
wire   [15:0] sub_ln703_267_fu_1872_p2;
wire   [15:0] add_ln703_399_fu_2342_p2;
wire   [15:0] add_ln703_398_fu_2337_p2;
wire   [15:0] sub_ln703_299_fu_2070_p2;
wire   [15:0] add_ln703_412_fu_2357_p2;
wire   [15:0] add_ln703_411_fu_2352_p2;
wire   [15:0] sub_ln703_315_fu_2188_p2;
wire   [15:0] add_ln703_414_fu_2367_p2;
wire   [15:0] sub_ln703_244_fu_1827_p2;
wire   [15:0] add_ln703_426_fu_2378_p2;
wire   [15:0] sub_ln703_313_fu_2413_p2;
wire   [15:0] sub_ln703_314_fu_2417_p2;
wire   [15:0] sub_ln703_316_fu_2421_p2;
wire   [15:0] add_ln703_368_fu_2429_p2;
wire   [15:0] add_ln703_370_fu_2437_p2;
wire   [15:0] sub_ln703_326_fu_2441_p2;
wire   [15:0] sub_ln703_312_fu_2409_p2;
wire   [15:0] add_ln703_373_fu_2445_p2;
wire   [15:0] sub_ln703_329_fu_2450_p2;
wire   [15:0] sub_ln703_317_fu_2425_p2;
wire   [15:0] sub_ln703_334_fu_2464_p2;
wire   [15:0] sub_ln703_336_fu_2469_p2;
wire   [15:0] sub_ln703_337_fu_2473_p2;
wire   [15:0] sub_ln703_338_fu_2478_p2;
wire   [15:0] sub_ln703_294_fu_2405_p2;
wire   [15:0] add_ln703_395_fu_2564_p2;
wire   [15:0] add_ln703_393_fu_2559_p2;
wire   [15:0] sub_ln703_339_fu_2482_p2;
wire   [15:0] add_ln703_382_fu_2486_p2;
wire   [15:0] add_ln703_383_fu_2490_p2;
wire   [15:0] sub_ln703_340_fu_2495_p2;
wire   [15:0] add_ln703_385_fu_2499_p2;
wire   [15:0] sub_ln703_341_fu_2504_p2;
wire   [15:0] sub_ln703_342_fu_2509_p2;
wire   [15:0] add_ln703_386_fu_2514_p2;
wire   [15:0] add_ln703_387_fu_2518_p2;
wire   [15:0] sub_ln703_344_fu_2523_p2;
wire   [15:0] add_ln703_391_fu_2527_p2;
wire   [15:0] sub_ln703_320_fu_2433_p2;
wire   [15:0] add_ln703_403_fu_2645_p2;
wire   [15:0] sub_ln703_347_fu_2536_p2;
wire   [15:0] add_ln703_392_fu_2540_p2;
wire   [15:0] sub_ln703_348_fu_2545_p2;
wire   [15:0] sub_ln703_350_fu_2554_p2;
wire   [15:0] add_ln703_407_fu_2675_p2;
wire   [15:0] add_ln703_396_fu_2568_p2;
wire   [15:0] sub_ln703_351_fu_2574_p2;
wire   [15:0] sub_ln703_352_fu_2579_p2;
wire   [15:0] sub_ln703_353_fu_2584_p2;
wire   [15:0] sub_ln703_354_fu_2589_p2;
wire   [15:0] sub_ln703_355_fu_2594_p2;
wire   [15:0] add_ln703_397_fu_2599_p2;
wire   [15:0] sub_ln703_358_fu_2613_p2;
wire   [15:0] sub_ln703_359_fu_2618_p2;
wire   [15:0] add_ln703_417_fu_2737_p2;
wire   [15:0] add_ln703_416_fu_2733_p2;
wire   [15:0] add_ln703_401_fu_2623_p2;
wire   [15:0] sub_ln703_360_fu_2627_p2;
wire   [15:0] add_ln703_419_fu_2757_p2;
wire   [15:0] sub_ln703_333_fu_2460_p2;
wire   [15:0] add_ln703_421_fu_2766_p2;
wire   [15:0] sub_ln703_362_fu_2641_p2;
wire   [15:0] add_ln703_405_fu_2650_p2;
wire   [15:0] add_ln703_406_fu_2655_p2;
wire   [15:0] sub_ln703_363_fu_2660_p2;
wire   [15:0] sub_ln703_364_fu_2665_p2;
wire   [15:0] add_ln703_408_fu_2679_p2;
wire   [15:0] sub_ln703_367_fu_2689_p2;
wire   [15:0] sub_ln703_368_fu_2694_p2;
wire   [15:0] add_ln703_409_fu_2704_p2;
wire   [15:0] add_ln703_429_fu_2825_p2;
wire   [15:0] add_ln703_430_fu_2829_p2;
wire   [15:0] sub_ln703_371_fu_2719_p2;
wire   [15:0] sub_ln703_373_fu_2723_p2;
wire   [15:0] sub_ln703_376_fu_2752_p2;
wire   [15:0] add_ln703_420_fu_2761_p2;
wire   [15:0] add_ln703_422_fu_2771_p2;
wire   [15:0] sub_ln703_378_fu_2776_p2;
wire   [15:0] sub_ln703_380_fu_2786_p2;
wire   [15:0] sub_ln703_382_fu_2796_p2;
wire   [15:0] sub_ln703_365_fu_2670_p2;
wire   [15:0] sub_ln703_370_fu_2714_p2;
wire   [15:0] sub_ln703_388_fu_2821_p2;
wire   [15:0] add_ln703_431_fu_2834_p2;
wire   [15:0] sub_ln703_391_fu_2844_p2;
wire   [15:0] sub_ln703_330_fu_2455_p2;
wire   [15:0] add_ln703_441_fu_2913_p2;
wire   [15:0] add_ln703_440_fu_2908_p2;
wire   [15:0] sub_ln703_396_fu_2858_p2;
wire   [15:0] sub_ln703_400_fu_2868_p2;
wire   [15:0] sub_ln703_383_fu_2801_p2;
wire   [15:0] add_ln703_438_fu_2888_p2;
wire   [15:0] sub_ln703_345_fu_2532_p2;
wire   [15:0] add_ln703_477_fu_2947_p2;
wire   [15:0] add_ln703_479_fu_2957_p2;
wire   [15:0] add_ln703_478_fu_2952_p2;
wire   [15:0] sub_ln703_395_fu_2853_p2;
wire   [15:0] sub_ln703_349_fu_2549_p2;
wire   [15:0] sub_ln703_372_fu_2985_p2;
wire   [15:0] sub_ln703_377_fu_2989_p2;
wire   [15:0] add_ln703_423_fu_2993_p2;
wire   [15:0] sub_ln703_384_fu_2997_p2;
wire   [15:0] add_ln703_425_fu_3001_p2;
wire   [15:0] sub_ln703_387_fu_3005_p2;
wire   [15:0] sub_ln703_390_fu_3009_p2;
wire   [15:0] add_ln703_432_fu_3014_p2;
wire   [15:0] sub_ln703_393_fu_3018_p2;
wire   [15:0] sub_ln703_394_fu_3022_p2;
wire   [15:0] sub_ln703_399_fu_3031_p2;
wire   [15:0] add_ln703_433_fu_3036_p2;
wire   [15:0] sub_ln703_401_fu_3040_p2;
wire   [15:0] sub_ln703_403_fu_3044_p2;
wire   [15:0] sub_ln703_404_fu_3049_p2;
wire   [15:0] add_ln703_437_fu_3053_p2;
wire   [15:0] sub_ln703_406_fu_3062_p2;
wire   [15:0] sub_ln703_410_fu_3071_p2;
wire   [15:0] add_ln703_439_fu_3075_p2;
wire   [15:0] add_ln703_450_fu_3168_p2;
wire   [15:0] sub_ln703_412_fu_3080_p2;
wire   [15:0] add_ln703_443_fu_3099_p2;
wire   [15:0] sub_ln703_417_fu_3103_p2;
wire   [15:0] sub_ln703_418_fu_3108_p2;
wire   [15:0] sub_ln703_419_fu_3113_p2;
wire   [15:0] sub_ln703_420_fu_3117_p2;
wire   [15:0] add_ln703_445_fu_3122_p2;
wire   [15:0] sub_ln703_424_fu_3140_p2;
wire   [15:0] add_ln703_455_fu_3237_p2;
wire   [15:0] sub_ln703_405_fu_3057_p2;
wire   [15:0] sub_ln703_425_fu_3145_p2;
wire   [15:0] add_ln703_448_fu_3150_p2;
wire   [15:0] sub_ln703_427_fu_3154_p2;
wire   [15:0] add_ln703_449_fu_3158_p2;
wire   [15:0] add_ln703_452_fu_3172_p2;
wire   [15:0] sub_ln703_429_fu_3177_p2;
wire   [15:0] sub_ln703_431_fu_3185_p2;
wire   [15:0] sub_ln703_413_fu_3084_p2;
wire   [15:0] sub_ln703_415_fu_3094_p2;
wire   [15:0] sub_ln703_432_fu_3190_p2;
wire   [15:0] sub_ln703_433_fu_3194_p2;
wire   [15:0] sub_ln703_436_fu_3208_p2;
wire   [15:0] sub_ln703_437_fu_3213_p2;
wire   [15:0] add_ln703_453_fu_3218_p2;
wire   [15:0] sub_ln703_438_fu_3223_p2;
wire   [15:0] sub_ln703_421_fu_3126_p2;
wire   [15:0] sub_ln703_439_fu_3228_p2;
wire   [15:0] sub_ln703_422_fu_3130_p2;
wire   [15:0] add_ln703_454_fu_3232_p2;
wire   [15:0] add_ln703_456_fu_3241_p2;
wire   [15:0] sub_ln703_440_fu_3247_p2;
wire   [15:0] sub_ln703_407_fu_3066_p2;
wire   [15:0] add_ln703_466_fu_3358_p2;
wire   [15:0] sub_ln703_441_fu_3252_p2;
wire   [15:0] sub_ln703_444_fu_3266_p2;
wire   [15:0] sub_ln703_445_fu_3271_p2;
wire   [15:0] sub_ln703_446_fu_3276_p2;
wire   [15:0] add_ln703_457_fu_3281_p2;
wire   [15:0] add_ln703_458_fu_3286_p2;
wire   [15:0] sub_ln703_414_fu_3089_p2;
wire   [15:0] add_ln703_470_fu_3398_p2;
wire   [15:0] add_ln703_459_fu_3292_p2;
wire   [15:0] sub_ln703_447_fu_3298_p2;
wire   [15:0] add_ln703_460_fu_3303_p2;
wire   [15:0] sub_ln703_398_fu_3026_p2;
wire   [15:0] add_ln703_474_fu_3428_p2;
wire   [15:0] add_ln703_473_fu_3423_p2;
wire   [15:0] add_ln703_461_fu_3323_p2;
wire   [15:0] sub_ln703_423_fu_3135_p2;
wire   [15:0] add_ln703_481_fu_3443_p2;
wire   [15:0] sub_ln703_442_fu_3256_p2;
wire   [15:0] sub_ln703_443_fu_3261_p2;
wire   [15:0] add_ln703_469_fu_3383_p2;
wire   [15:0] sub_ln703_430_fu_3181_p2;
wire   [15:0] add_ln703_489_fu_3468_p2;
wire   [15:0] add_ln703_472_fu_3413_p2;
wire   [15:0] sub_ln703_435_fu_3204_p2;
wire   [15:0] add_ln703_494_fu_3487_p2;
wire   [15:0] sub_ln703_449_fu_3313_p2;
wire   [15:0] add_ln703_486_fu_3453_p2;
wire   [15:0] add_ln703_487_fu_3458_p2;
wire   [15:0] add_ln703_490_fu_3473_p2;
wire   [15:0] add_ln703_495_fu_3492_p2;
wire   [15:0] add_ln703_476_fu_3531_p2;
wire   [15:0] sub_ln703_460_fu_3535_p2;
wire   [15:0] sub_ln703_462_fu_3539_p2;
wire   [15:0] sub_ln703_463_fu_3543_p2;
wire   [15:0] sub_ln703_464_fu_3547_p2;
wire   [15:0] sub_ln703_465_fu_3551_p2;
wire   [15:0] add_ln703_484_fu_3555_p2;
wire   [15:0] add_ln703_485_fu_3559_p2;
wire   [15:0] sub_ln703_466_fu_3563_p2;
wire   [15:0] sub_ln703_467_fu_3567_p2;
wire   [15:0] add_ln703_488_fu_3571_p2;
wire   [15:0] sub_ln703_468_fu_3575_p2;
wire   [15:0] sub_ln703_470_fu_3579_p2;
wire   [15:0] sub_ln703_471_fu_3583_p2;
wire   [15:0] sub_ln703_472_fu_3587_p2;
wire   [15:0] sub_ln703_473_fu_3591_p2;
wire   [15:0] add_ln703_493_fu_3595_p2;
wire   [15:0] sub_ln703_475_fu_3599_p2;
wire   [15:0] sub_ln703_476_fu_3603_p2;
wire   [15:0] sub_ln703_477_fu_3607_p2;
wire   [15:0] sub_ln703_478_fu_3612_p2;
wire   [15:0] add_ln703_498_fu_3616_p2;
wire   [15:0] sub_ln703_479_fu_3621_p2;
wire   [15:0] sub_ln703_480_fu_3626_p2;
wire   [15:0] add_ln703_499_fu_3631_p2;
wire   [15:0] sub_ln703_482_fu_3640_p2;
wire   [15:0] sub_ln703_483_fu_3645_p2;
wire   [15:0] sub_ln703_484_fu_3650_p2;
wire   [15:0] add_ln703_500_fu_3655_p2;
wire   [15:0] sub_ln703_485_fu_3660_p2;
wire   [15:0] sub_ln703_488_fu_3665_p2;
wire   [15:0] sub_ln703_489_fu_3670_p2;
wire   [15:0] sub_ln703_492_fu_3679_p2;
wire   [15:0] sub_ln703_493_fu_3684_p2;
wire   [15:0] sub_ln703_494_fu_3689_p2;
wire   [15:0] sub_ln703_495_fu_3694_p2;
wire   [15:0] sub_ln703_496_fu_3699_p2;
wire   [15:0] add_ln703_501_fu_3708_p2;
wire   [15:0] add_ln703_502_fu_3713_p2;
wire   [15:0] sub_ln703_499_fu_3723_p2;
wire   [15:0] add_ln703_508_fu_3843_p2;
wire   [15:0] sub_ln703_501_fu_3728_p2;
wire   [15:0] sub_ln703_502_fu_3732_p2;
wire   [15:0] add_ln703_514_fu_3862_p2;
wire   [15:0] add_ln703_518_fu_3875_p2;
wire   [15:0] add_ln703_517_fu_3871_p2;
wire   [15:0] sub_ln703_503_fu_3737_p2;
wire   [15:0] sub_ln703_504_fu_3742_p2;
wire   [15:0] sub_ln703_505_fu_3747_p2;
wire   [15:0] sub_ln703_481_fu_3636_p2;
wire   [15:0] sub_ln703_506_fu_3752_p2;
wire   [15:0] add_ln703_503_fu_3757_p2;
wire   [15:0] sub_ln703_507_fu_3762_p2;
wire   [15:0] sub_ln703_508_fu_3767_p2;
wire   [15:0] sub_ln703_509_fu_3772_p2;
wire   [15:0] add_ln703_504_fu_3777_p2;
wire   [15:0] sub_ln703_510_fu_3781_p2;
wire   [15:0] add_ln703_505_fu_3785_p2;
wire   [15:0] add_ln703_527_fu_3949_p2;
wire   [15:0] add_ln703_526_fu_3945_p2;
wire   [15:0] sub_ln703_511_fu_3790_p2;
wire   [15:0] sub_ln703_490_fu_3675_p2;
wire   [15:0] add_ln703_506_fu_3795_p2;
wire   [15:0] add_ln703_507_fu_3799_p2;
wire   [15:0] sub_ln703_512_fu_3804_p2;
wire   [15:0] sub_ln703_513_fu_3809_p2;
wire   [15:0] sub_ln703_514_fu_3814_p2;
wire   [15:0] sub_ln703_515_fu_3819_p2;
wire   [15:0] sub_ln703_497_fu_3704_p2;
wire   [15:0] sub_ln703_516_fu_3824_p2;
wire   [15:0] sub_ln703_517_fu_3829_p2;
wire   [15:0] sub_ln703_498_fu_3718_p2;
wire   [15:0] sub_ln703_518_fu_3834_p2;
wire   [15:0] sub_ln703_519_fu_3839_p2;
wire   [15:0] add_ln703_511_fu_3847_p2;
wire   [15:0] acc_1_V_fu_3852_p2;
wire   [15:0] acc_2_V_fu_3857_p2;
wire   [15:0] acc_3_V_fu_3866_p2;
wire   [15:0] acc_4_V_fu_3879_p2;
wire   [15:0] acc_5_V_fu_3885_p2;
wire   [15:0] acc_6_V_fu_3890_p2;
wire   [15:0] acc_7_V_fu_3895_p2;
wire   [15:0] acc_8_V_fu_3900_p2;
wire   [15:0] acc_9_V_fu_3905_p2;
wire   [15:0] acc_10_V_fu_3910_p2;
wire   [15:0] acc_11_V_fu_3915_p2;
wire   [15:0] acc_12_V_fu_3920_p2;
wire   [15:0] acc_13_V_fu_3925_p2;
wire   [15:0] acc_14_V_fu_3930_p2;
wire   [15:0] acc_15_V_fu_3935_p2;
wire   [15:0] acc_16_V_fu_3940_p2;
wire   [15:0] acc_17_V_fu_3953_p2;
wire   [15:0] acc_18_V_fu_3959_p2;
wire   [15:0] acc_19_V_fu_3964_p2;
wire   [15:0] acc_20_V_fu_3969_p2;
wire   [15:0] acc_21_V_fu_3974_p2;
wire   [15:0] acc_22_V_fu_3979_p2;
wire   [15:0] acc_23_V_fu_3984_p2;
wire   [15:0] acc_24_V_fu_3989_p2;
wire   [15:0] acc_25_V_fu_3994_p2;
wire   [15:0] acc_26_V_fu_3999_p2;
wire   [15:0] acc_27_V_fu_4004_p2;
wire   [15:0] acc_28_V_fu_4009_p2;
wire   [15:0] acc_29_V_fu_4014_p2;
wire   [15:0] acc_30_V_fu_4019_p2;
wire   [15:0] acc_31_V_fu_4024_p2;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        add_ln703_200_reg_5077 <= add_ln703_200_fu_304_p2;
        add_ln703_200_reg_5077_pp0_iter2_reg <= add_ln703_200_reg_5077;
        add_ln703_201_reg_5090 <= add_ln703_201_fu_312_p2;
        add_ln703_201_reg_5090_pp0_iter2_reg <= add_ln703_201_reg_5090;
        add_ln703_202_reg_5096 <= add_ln703_202_fu_316_p2;
        add_ln703_202_reg_5096_pp0_iter2_reg <= add_ln703_202_reg_5096;
        add_ln703_203_reg_5113 <= add_ln703_203_fu_329_p2;
        add_ln703_204_reg_5101 <= add_ln703_204_fu_320_p2;
        add_ln703_204_reg_5101_pp0_iter2_reg <= add_ln703_204_reg_5101;
        add_ln703_205_reg_5119 <= add_ln703_205_fu_333_p2;
        add_ln703_206_reg_5131 <= add_ln703_206_fu_341_p2;
        add_ln703_207_reg_5107 <= add_ln703_207_fu_325_p2;
        add_ln703_207_reg_5107_pp0_iter2_reg <= add_ln703_207_reg_5107;
        add_ln703_208_reg_5137 <= add_ln703_208_fu_345_p2;
        add_ln703_209_reg_5178 <= add_ln703_209_fu_416_p2;
        add_ln703_210_reg_5143 <= add_ln703_210_fu_349_p2;
        add_ln703_210_reg_5143_pp0_iter3_reg <= add_ln703_210_reg_5143;
        add_ln703_211_reg_5184 <= add_ln703_211_fu_420_p2;
        add_ln703_213_reg_5189 <= add_ln703_213_fu_429_p2;
        add_ln703_214_reg_5194 <= add_ln703_214_fu_433_p2;
        add_ln703_216_reg_5215 <= add_ln703_216_fu_461_p2;
        add_ln703_220_reg_5221 <= add_ln703_220_fu_484_p2;
        add_ln703_223_reg_5231 <= add_ln703_223_fu_507_p2;
        add_ln703_225_reg_5237 <= add_ln703_225_fu_513_p2;
        add_ln703_227_reg_5242 <= add_ln703_227_fu_522_p2;
        add_ln703_233_reg_5149 <= add_ln703_233_fu_353_p2;
        add_ln703_233_reg_5149_pp0_iter3_reg <= add_ln703_233_reg_5149;
        add_ln703_234_reg_5264 <= add_ln703_234_fu_564_p2;
        add_ln703_238_reg_5269 <= add_ln703_238_fu_569_p2;
        add_ln703_246_reg_5320 <= add_ln703_246_fu_787_p2;
        add_ln703_247_reg_5159 <= add_ln703_247_fu_357_p2;
        add_ln703_247_reg_5159_pp0_iter3_reg <= add_ln703_247_reg_5159;
        add_ln703_251_reg_5289 <= add_ln703_251_fu_589_p2;
        add_ln703_258_reg_5295 <= add_ln703_258_fu_593_p2;
        add_ln703_261_reg_5360 <= add_ln703_261_fu_955_p2;
        add_ln703_267_reg_5405 <= add_ln703_267_fu_1055_p2;
        add_ln703_268_reg_5415 <= add_ln703_268_fu_1065_p2;
        add_ln703_272_reg_5304 <= add_ln703_272_fu_597_p2;
        add_ln703_272_reg_5304_pp0_iter4_reg <= add_ln703_272_reg_5304;
        add_ln703_274_reg_5420 <= add_ln703_274_fu_1089_p2;
        add_ln703_276_reg_5430 <= add_ln703_276_fu_1100_p2;
        add_ln703_278_reg_5435 <= add_ln703_278_fu_1105_p2;
        add_ln703_281_reg_5455 <= add_ln703_281_fu_1129_p2;
        add_ln703_283_reg_5460 <= add_ln703_283_fu_1140_p2;
        add_ln703_287_reg_5525 <= add_ln703_287_fu_1354_p2;
        add_ln703_288_reg_5475 <= add_ln703_288_fu_1156_p2;
        add_ln703_291_reg_5530 <= add_ln703_291_fu_1371_p2;
        add_ln703_301_reg_5550 <= add_ln703_301_fu_1494_p2;
        add_ln703_304_reg_5314 <= add_ln703_304_fu_601_p2;
        add_ln703_307_reg_5555 <= add_ln703_307_fu_1504_p2;
        add_ln703_309_reg_5484 <= add_ln703_309_fu_1179_p2;
        add_ln703_314_reg_5490 <= add_ln703_314_fu_1183_p2;
        add_ln703_316_reg_5496 <= add_ln703_316_fu_1187_p2;
        add_ln703_321_reg_5590 <= add_ln703_321_fu_1636_p2;
        add_ln703_323_reg_5506 <= add_ln703_323_fu_1198_p2;
        add_ln703_326_reg_5625 <= add_ln703_326_fu_1686_p2;
        add_ln703_330_reg_5640 <= add_ln703_330_fu_1710_p2;
        add_ln703_335_reg_5645 <= add_ln703_335_fu_1730_p2;
        add_ln703_339_reg_5655 <= add_ln703_339_fu_1740_p2;
        add_ln703_343_reg_5660 <= add_ln703_343_fu_1745_p2;
        add_ln703_347_reg_5675 <= add_ln703_347_fu_1760_p2;
        add_ln703_353_reg_5743 <= add_ln703_353_fu_2060_p2;
        add_ln703_354_reg_5753 <= add_ln703_354_fu_2080_p2;
        add_ln703_357_reg_5683 <= add_ln703_357_fu_1764_p2;
        add_ln703_357_reg_5683_pp0_iter6_reg <= add_ln703_357_reg_5683;
        add_ln703_359_reg_5768 <= add_ln703_359_fu_2127_p2;
        add_ln703_371_reg_5691 <= add_ln703_371_fu_1768_p2;
        add_ln703_372_reg_5793 <= add_ln703_372_fu_2228_p2;
        add_ln703_377_reg_5833 <= add_ln703_377_fu_2283_p2;
        add_ln703_379_reg_5838 <= add_ln703_379_fu_2292_p2;
        add_ln703_381_reg_5848 <= add_ln703_381_fu_2307_p2;
        add_ln703_384_reg_5701 <= add_ln703_384_fu_1772_p2;
        add_ln703_384_reg_5701_pp0_iter6_reg <= add_ln703_384_reg_5701;
        add_ln703_390_reg_5858 <= add_ln703_390_fu_2326_p2;
        add_ln703_394_reg_5710 <= add_ln703_394_fu_1776_p2;
        add_ln703_394_reg_5710_pp0_iter6_reg <= add_ln703_394_reg_5710;
        add_ln703_400_reg_5868 <= add_ln703_400_fu_2346_p2;
        add_ln703_402_reg_5931 <= add_ln703_402_fu_2631_p2;
        add_ln703_404_reg_5718 <= add_ln703_404_fu_1780_p2;
        add_ln703_404_reg_5718_pp0_iter6_reg <= add_ln703_404_reg_5718;
        add_ln703_410_reg_5951 <= add_ln703_410_fu_2709_p2;
        add_ln703_413_reg_5873 <= add_ln703_413_fu_2361_p2;
        add_ln703_415_reg_5878 <= add_ln703_415_fu_2372_p2;
        add_ln703_418_reg_5961 <= add_ln703_418_fu_2741_p2;
        add_ln703_424_reg_5981 <= add_ln703_424_fu_2806_p2;
        add_ln703_427_reg_5883 <= add_ln703_427_fu_2383_p2;
        add_ln703_428_reg_5888 <= add_ln703_428_fu_2389_p2;
        add_ln703_434_reg_6011 <= add_ln703_434_fu_2873_p2;
        add_ln703_435_reg_5894 <= add_ln703_435_fu_2393_p2;
        add_ln703_436_reg_6021 <= add_ln703_436_fu_2883_p2;
        add_ln703_442_reg_6041 <= add_ln703_442_fu_2917_p2;
        add_ln703_444_reg_6051 <= add_ln703_444_fu_2928_p2;
        add_ln703_446_reg_5901 <= add_ln703_446_fu_2397_p2;
        add_ln703_447_reg_6056 <= add_ln703_447_fu_2933_p2;
        add_ln703_451_reg_6066 <= add_ln703_451_fu_2943_p2;
        add_ln703_451_reg_6066_pp0_iter8_reg <= add_ln703_451_reg_6066;
        add_ln703_462_reg_5909 <= add_ln703_462_fu_2401_p2;
        add_ln703_462_reg_5909_pp0_iter7_reg <= add_ln703_462_reg_5909;
        add_ln703_462_reg_5909_pp0_iter8_reg <= add_ln703_462_reg_5909_pp0_iter7_reg;
        add_ln703_463_reg_6128 <= add_ln703_463_fu_3328_p2;
        add_ln703_464_reg_6133 <= add_ln703_464_fu_3333_p2;
        add_ln703_465_reg_6138 <= add_ln703_465_fu_3338_p2;
        add_ln703_467_reg_6158 <= add_ln703_467_fu_3363_p2;
        add_ln703_468_reg_6173 <= add_ln703_468_fu_3378_p2;
        add_ln703_471_reg_6188 <= add_ln703_471_fu_3403_p2;
        add_ln703_475_reg_6203 <= add_ln703_475_fu_3432_p2;
        add_ln703_480_reg_6072 <= add_ln703_480_fu_2961_p2;
        add_ln703_480_reg_6072_pp0_iter8_reg <= add_ln703_480_reg_6072;
        add_ln703_482_reg_6077 <= add_ln703_482_fu_2967_p2;
        add_ln703_483_reg_6213 <= add_ln703_483_fu_3448_p2;
        add_ln703_491_reg_6087 <= add_ln703_491_fu_2971_p2;
        add_ln703_491_reg_6087_pp0_iter8_reg <= add_ln703_491_reg_6087;
        add_ln703_492_reg_6223 <= add_ln703_492_fu_3478_p2;
        add_ln703_496_reg_6234 <= add_ln703_496_fu_3497_p2;
        add_ln703_497_reg_6239 <= add_ln703_497_fu_3501_p2;
        add_ln703_509_reg_6092 <= add_ln703_509_fu_2976_p2;
        add_ln703_509_reg_6092_pp0_iter8_reg <= add_ln703_509_reg_6092;
        add_ln703_510_reg_6264 <= add_ln703_510_fu_3527_p2;
        add_ln703_516_reg_6103 <= add_ln703_516_fu_2980_p2;
        add_ln703_516_reg_6103_pp0_iter8_reg <= add_ln703_516_reg_6103;
        add_ln703_reg_5052 <= add_ln703_fu_280_p2;
        data_10_V_read11_reg_4832 <= data_10_V_read_int_reg;
        data_10_V_read11_reg_4832_pp0_iter1_reg <= data_10_V_read11_reg_4832;
        data_10_V_read11_reg_4832_pp0_iter2_reg <= data_10_V_read11_reg_4832_pp0_iter1_reg;
        data_10_V_read11_reg_4832_pp0_iter3_reg <= data_10_V_read11_reg_4832_pp0_iter2_reg;
        data_10_V_read11_reg_4832_pp0_iter4_reg <= data_10_V_read11_reg_4832_pp0_iter3_reg;
        data_11_V_read12_reg_4808 <= data_11_V_read_int_reg;
        data_11_V_read12_reg_4808_pp0_iter1_reg <= data_11_V_read12_reg_4808;
        data_11_V_read12_reg_4808_pp0_iter2_reg <= data_11_V_read12_reg_4808_pp0_iter1_reg;
        data_11_V_read12_reg_4808_pp0_iter3_reg <= data_11_V_read12_reg_4808_pp0_iter2_reg;
        data_11_V_read12_reg_4808_pp0_iter4_reg <= data_11_V_read12_reg_4808_pp0_iter3_reg;
        data_12_V_read13_reg_4778 <= data_12_V_read_int_reg;
        data_12_V_read13_reg_4778_pp0_iter1_reg <= data_12_V_read13_reg_4778;
        data_12_V_read13_reg_4778_pp0_iter2_reg <= data_12_V_read13_reg_4778_pp0_iter1_reg;
        data_12_V_read13_reg_4778_pp0_iter3_reg <= data_12_V_read13_reg_4778_pp0_iter2_reg;
        data_12_V_read13_reg_4778_pp0_iter4_reg <= data_12_V_read13_reg_4778_pp0_iter3_reg;
        data_13_V_read14_reg_4745 <= data_13_V_read_int_reg;
        data_13_V_read14_reg_4745_pp0_iter1_reg <= data_13_V_read14_reg_4745;
        data_13_V_read14_reg_4745_pp0_iter2_reg <= data_13_V_read14_reg_4745_pp0_iter1_reg;
        data_13_V_read14_reg_4745_pp0_iter3_reg <= data_13_V_read14_reg_4745_pp0_iter2_reg;
        data_13_V_read14_reg_4745_pp0_iter4_reg <= data_13_V_read14_reg_4745_pp0_iter3_reg;
        data_13_V_read14_reg_4745_pp0_iter5_reg <= data_13_V_read14_reg_4745_pp0_iter4_reg;
        data_14_V_read15_reg_4714 <= data_14_V_read_int_reg;
        data_14_V_read15_reg_4714_pp0_iter1_reg <= data_14_V_read15_reg_4714;
        data_14_V_read15_reg_4714_pp0_iter2_reg <= data_14_V_read15_reg_4714_pp0_iter1_reg;
        data_14_V_read15_reg_4714_pp0_iter3_reg <= data_14_V_read15_reg_4714_pp0_iter2_reg;
        data_14_V_read15_reg_4714_pp0_iter4_reg <= data_14_V_read15_reg_4714_pp0_iter3_reg;
        data_14_V_read15_reg_4714_pp0_iter5_reg <= data_14_V_read15_reg_4714_pp0_iter4_reg;
        data_15_V_read16_reg_4682 <= data_15_V_read_int_reg;
        data_15_V_read16_reg_4682_pp0_iter1_reg <= data_15_V_read16_reg_4682;
        data_15_V_read16_reg_4682_pp0_iter2_reg <= data_15_V_read16_reg_4682_pp0_iter1_reg;
        data_15_V_read16_reg_4682_pp0_iter3_reg <= data_15_V_read16_reg_4682_pp0_iter2_reg;
        data_15_V_read16_reg_4682_pp0_iter4_reg <= data_15_V_read16_reg_4682_pp0_iter3_reg;
        data_15_V_read16_reg_4682_pp0_iter5_reg <= data_15_V_read16_reg_4682_pp0_iter4_reg;
        data_16_V_read17_reg_4650 <= data_16_V_read_int_reg;
        data_16_V_read17_reg_4650_pp0_iter1_reg <= data_16_V_read17_reg_4650;
        data_16_V_read17_reg_4650_pp0_iter2_reg <= data_16_V_read17_reg_4650_pp0_iter1_reg;
        data_16_V_read17_reg_4650_pp0_iter3_reg <= data_16_V_read17_reg_4650_pp0_iter2_reg;
        data_16_V_read17_reg_4650_pp0_iter4_reg <= data_16_V_read17_reg_4650_pp0_iter3_reg;
        data_16_V_read17_reg_4650_pp0_iter5_reg <= data_16_V_read17_reg_4650_pp0_iter4_reg;
        data_17_V_read_8_reg_4621 <= data_17_V_read_int_reg;
        data_17_V_read_8_reg_4621_pp0_iter1_reg <= data_17_V_read_8_reg_4621;
        data_17_V_read_8_reg_4621_pp0_iter2_reg <= data_17_V_read_8_reg_4621_pp0_iter1_reg;
        data_17_V_read_8_reg_4621_pp0_iter3_reg <= data_17_V_read_8_reg_4621_pp0_iter2_reg;
        data_17_V_read_8_reg_4621_pp0_iter4_reg <= data_17_V_read_8_reg_4621_pp0_iter3_reg;
        data_17_V_read_8_reg_4621_pp0_iter5_reg <= data_17_V_read_8_reg_4621_pp0_iter4_reg;
        data_17_V_read_8_reg_4621_pp0_iter6_reg <= data_17_V_read_8_reg_4621_pp0_iter5_reg;
        data_18_V_read_7_reg_4594 <= data_18_V_read_int_reg;
        data_18_V_read_7_reg_4594_pp0_iter1_reg <= data_18_V_read_7_reg_4594;
        data_18_V_read_7_reg_4594_pp0_iter2_reg <= data_18_V_read_7_reg_4594_pp0_iter1_reg;
        data_18_V_read_7_reg_4594_pp0_iter3_reg <= data_18_V_read_7_reg_4594_pp0_iter2_reg;
        data_18_V_read_7_reg_4594_pp0_iter4_reg <= data_18_V_read_7_reg_4594_pp0_iter3_reg;
        data_18_V_read_7_reg_4594_pp0_iter5_reg <= data_18_V_read_7_reg_4594_pp0_iter4_reg;
        data_18_V_read_7_reg_4594_pp0_iter6_reg <= data_18_V_read_7_reg_4594_pp0_iter5_reg;
        data_19_V_read_7_reg_4567 <= data_19_V_read_int_reg;
        data_19_V_read_7_reg_4567_pp0_iter1_reg <= data_19_V_read_7_reg_4567;
        data_19_V_read_7_reg_4567_pp0_iter2_reg <= data_19_V_read_7_reg_4567_pp0_iter1_reg;
        data_19_V_read_7_reg_4567_pp0_iter3_reg <= data_19_V_read_7_reg_4567_pp0_iter2_reg;
        data_19_V_read_7_reg_4567_pp0_iter4_reg <= data_19_V_read_7_reg_4567_pp0_iter3_reg;
        data_19_V_read_7_reg_4567_pp0_iter5_reg <= data_19_V_read_7_reg_4567_pp0_iter4_reg;
        data_19_V_read_7_reg_4567_pp0_iter6_reg <= data_19_V_read_7_reg_4567_pp0_iter5_reg;
        data_20_V_read21_reg_4539 <= data_20_V_read_int_reg;
        data_20_V_read21_reg_4539_pp0_iter1_reg <= data_20_V_read21_reg_4539;
        data_20_V_read21_reg_4539_pp0_iter2_reg <= data_20_V_read21_reg_4539_pp0_iter1_reg;
        data_20_V_read21_reg_4539_pp0_iter3_reg <= data_20_V_read21_reg_4539_pp0_iter2_reg;
        data_20_V_read21_reg_4539_pp0_iter4_reg <= data_20_V_read21_reg_4539_pp0_iter3_reg;
        data_20_V_read21_reg_4539_pp0_iter5_reg <= data_20_V_read21_reg_4539_pp0_iter4_reg;
        data_20_V_read21_reg_4539_pp0_iter6_reg <= data_20_V_read21_reg_4539_pp0_iter5_reg;
        data_21_V_read22_reg_4512 <= data_21_V_read_int_reg;
        data_21_V_read22_reg_4512_pp0_iter1_reg <= data_21_V_read22_reg_4512;
        data_21_V_read22_reg_4512_pp0_iter2_reg <= data_21_V_read22_reg_4512_pp0_iter1_reg;
        data_21_V_read22_reg_4512_pp0_iter3_reg <= data_21_V_read22_reg_4512_pp0_iter2_reg;
        data_21_V_read22_reg_4512_pp0_iter4_reg <= data_21_V_read22_reg_4512_pp0_iter3_reg;
        data_21_V_read22_reg_4512_pp0_iter5_reg <= data_21_V_read22_reg_4512_pp0_iter4_reg;
        data_21_V_read22_reg_4512_pp0_iter6_reg <= data_21_V_read22_reg_4512_pp0_iter5_reg;
        data_22_V_read23_reg_4483 <= data_22_V_read_int_reg;
        data_22_V_read23_reg_4483_pp0_iter1_reg <= data_22_V_read23_reg_4483;
        data_22_V_read23_reg_4483_pp0_iter2_reg <= data_22_V_read23_reg_4483_pp0_iter1_reg;
        data_22_V_read23_reg_4483_pp0_iter3_reg <= data_22_V_read23_reg_4483_pp0_iter2_reg;
        data_22_V_read23_reg_4483_pp0_iter4_reg <= data_22_V_read23_reg_4483_pp0_iter3_reg;
        data_22_V_read23_reg_4483_pp0_iter5_reg <= data_22_V_read23_reg_4483_pp0_iter4_reg;
        data_22_V_read23_reg_4483_pp0_iter6_reg <= data_22_V_read23_reg_4483_pp0_iter5_reg;
        data_22_V_read23_reg_4483_pp0_iter7_reg <= data_22_V_read23_reg_4483_pp0_iter6_reg;
        data_23_V_read24_reg_4451 <= data_23_V_read_int_reg;
        data_23_V_read24_reg_4451_pp0_iter1_reg <= data_23_V_read24_reg_4451;
        data_23_V_read24_reg_4451_pp0_iter2_reg <= data_23_V_read24_reg_4451_pp0_iter1_reg;
        data_23_V_read24_reg_4451_pp0_iter3_reg <= data_23_V_read24_reg_4451_pp0_iter2_reg;
        data_23_V_read24_reg_4451_pp0_iter4_reg <= data_23_V_read24_reg_4451_pp0_iter3_reg;
        data_23_V_read24_reg_4451_pp0_iter5_reg <= data_23_V_read24_reg_4451_pp0_iter4_reg;
        data_23_V_read24_reg_4451_pp0_iter6_reg <= data_23_V_read24_reg_4451_pp0_iter5_reg;
        data_23_V_read24_reg_4451_pp0_iter7_reg <= data_23_V_read24_reg_4451_pp0_iter6_reg;
        data_24_V_read25_reg_4421 <= data_24_V_read_int_reg;
        data_24_V_read25_reg_4421_pp0_iter1_reg <= data_24_V_read25_reg_4421;
        data_24_V_read25_reg_4421_pp0_iter2_reg <= data_24_V_read25_reg_4421_pp0_iter1_reg;
        data_24_V_read25_reg_4421_pp0_iter3_reg <= data_24_V_read25_reg_4421_pp0_iter2_reg;
        data_24_V_read25_reg_4421_pp0_iter4_reg <= data_24_V_read25_reg_4421_pp0_iter3_reg;
        data_24_V_read25_reg_4421_pp0_iter5_reg <= data_24_V_read25_reg_4421_pp0_iter4_reg;
        data_24_V_read25_reg_4421_pp0_iter6_reg <= data_24_V_read25_reg_4421_pp0_iter5_reg;
        data_24_V_read25_reg_4421_pp0_iter7_reg <= data_24_V_read25_reg_4421_pp0_iter6_reg;
        data_25_V_read26_reg_4391 <= data_25_V_read_int_reg;
        data_25_V_read26_reg_4391_pp0_iter1_reg <= data_25_V_read26_reg_4391;
        data_25_V_read26_reg_4391_pp0_iter2_reg <= data_25_V_read26_reg_4391_pp0_iter1_reg;
        data_25_V_read26_reg_4391_pp0_iter3_reg <= data_25_V_read26_reg_4391_pp0_iter2_reg;
        data_25_V_read26_reg_4391_pp0_iter4_reg <= data_25_V_read26_reg_4391_pp0_iter3_reg;
        data_25_V_read26_reg_4391_pp0_iter5_reg <= data_25_V_read26_reg_4391_pp0_iter4_reg;
        data_25_V_read26_reg_4391_pp0_iter6_reg <= data_25_V_read26_reg_4391_pp0_iter5_reg;
        data_25_V_read26_reg_4391_pp0_iter7_reg <= data_25_V_read26_reg_4391_pp0_iter6_reg;
        data_26_V_read27_reg_4365 <= data_26_V_read_int_reg;
        data_26_V_read27_reg_4365_pp0_iter1_reg <= data_26_V_read27_reg_4365;
        data_26_V_read27_reg_4365_pp0_iter2_reg <= data_26_V_read27_reg_4365_pp0_iter1_reg;
        data_26_V_read27_reg_4365_pp0_iter3_reg <= data_26_V_read27_reg_4365_pp0_iter2_reg;
        data_26_V_read27_reg_4365_pp0_iter4_reg <= data_26_V_read27_reg_4365_pp0_iter3_reg;
        data_26_V_read27_reg_4365_pp0_iter5_reg <= data_26_V_read27_reg_4365_pp0_iter4_reg;
        data_26_V_read27_reg_4365_pp0_iter6_reg <= data_26_V_read27_reg_4365_pp0_iter5_reg;
        data_26_V_read27_reg_4365_pp0_iter7_reg <= data_26_V_read27_reg_4365_pp0_iter6_reg;
        data_27_V_read_8_reg_4342 <= data_27_V_read_int_reg;
        data_27_V_read_8_reg_4342_pp0_iter1_reg <= data_27_V_read_8_reg_4342;
        data_27_V_read_8_reg_4342_pp0_iter2_reg <= data_27_V_read_8_reg_4342_pp0_iter1_reg;
        data_27_V_read_8_reg_4342_pp0_iter3_reg <= data_27_V_read_8_reg_4342_pp0_iter2_reg;
        data_27_V_read_8_reg_4342_pp0_iter4_reg <= data_27_V_read_8_reg_4342_pp0_iter3_reg;
        data_27_V_read_8_reg_4342_pp0_iter5_reg <= data_27_V_read_8_reg_4342_pp0_iter4_reg;
        data_27_V_read_8_reg_4342_pp0_iter6_reg <= data_27_V_read_8_reg_4342_pp0_iter5_reg;
        data_27_V_read_8_reg_4342_pp0_iter7_reg <= data_27_V_read_8_reg_4342_pp0_iter6_reg;
        data_28_V_read_7_reg_4313 <= data_28_V_read_int_reg;
        data_28_V_read_7_reg_4313_pp0_iter1_reg <= data_28_V_read_7_reg_4313;
        data_28_V_read_7_reg_4313_pp0_iter2_reg <= data_28_V_read_7_reg_4313_pp0_iter1_reg;
        data_28_V_read_7_reg_4313_pp0_iter3_reg <= data_28_V_read_7_reg_4313_pp0_iter2_reg;
        data_28_V_read_7_reg_4313_pp0_iter4_reg <= data_28_V_read_7_reg_4313_pp0_iter3_reg;
        data_28_V_read_7_reg_4313_pp0_iter5_reg <= data_28_V_read_7_reg_4313_pp0_iter4_reg;
        data_28_V_read_7_reg_4313_pp0_iter6_reg <= data_28_V_read_7_reg_4313_pp0_iter5_reg;
        data_28_V_read_7_reg_4313_pp0_iter7_reg <= data_28_V_read_7_reg_4313_pp0_iter6_reg;
        data_28_V_read_7_reg_4313_pp0_iter8_reg <= data_28_V_read_7_reg_4313_pp0_iter7_reg;
        data_29_V_read_7_reg_4279 <= data_29_V_read_int_reg;
        data_29_V_read_7_reg_4279_pp0_iter1_reg <= data_29_V_read_7_reg_4279;
        data_29_V_read_7_reg_4279_pp0_iter2_reg <= data_29_V_read_7_reg_4279_pp0_iter1_reg;
        data_29_V_read_7_reg_4279_pp0_iter3_reg <= data_29_V_read_7_reg_4279_pp0_iter2_reg;
        data_29_V_read_7_reg_4279_pp0_iter4_reg <= data_29_V_read_7_reg_4279_pp0_iter3_reg;
        data_29_V_read_7_reg_4279_pp0_iter5_reg <= data_29_V_read_7_reg_4279_pp0_iter4_reg;
        data_29_V_read_7_reg_4279_pp0_iter6_reg <= data_29_V_read_7_reg_4279_pp0_iter5_reg;
        data_29_V_read_7_reg_4279_pp0_iter7_reg <= data_29_V_read_7_reg_4279_pp0_iter6_reg;
        data_29_V_read_7_reg_4279_pp0_iter8_reg <= data_29_V_read_7_reg_4279_pp0_iter7_reg;
        data_2_V_read_9_reg_5035 <= data_2_V_read_int_reg;
        data_30_V_read31_reg_4250 <= data_30_V_read_int_reg;
        data_30_V_read31_reg_4250_pp0_iter1_reg <= data_30_V_read31_reg_4250;
        data_30_V_read31_reg_4250_pp0_iter2_reg <= data_30_V_read31_reg_4250_pp0_iter1_reg;
        data_30_V_read31_reg_4250_pp0_iter3_reg <= data_30_V_read31_reg_4250_pp0_iter2_reg;
        data_30_V_read31_reg_4250_pp0_iter4_reg <= data_30_V_read31_reg_4250_pp0_iter3_reg;
        data_30_V_read31_reg_4250_pp0_iter5_reg <= data_30_V_read31_reg_4250_pp0_iter4_reg;
        data_30_V_read31_reg_4250_pp0_iter6_reg <= data_30_V_read31_reg_4250_pp0_iter5_reg;
        data_30_V_read31_reg_4250_pp0_iter7_reg <= data_30_V_read31_reg_4250_pp0_iter6_reg;
        data_30_V_read31_reg_4250_pp0_iter8_reg <= data_30_V_read31_reg_4250_pp0_iter7_reg;
        data_31_V_read32_reg_4221 <= data_31_V_read_int_reg;
        data_31_V_read32_reg_4221_pp0_iter1_reg <= data_31_V_read32_reg_4221;
        data_31_V_read32_reg_4221_pp0_iter2_reg <= data_31_V_read32_reg_4221_pp0_iter1_reg;
        data_31_V_read32_reg_4221_pp0_iter3_reg <= data_31_V_read32_reg_4221_pp0_iter2_reg;
        data_31_V_read32_reg_4221_pp0_iter4_reg <= data_31_V_read32_reg_4221_pp0_iter3_reg;
        data_31_V_read32_reg_4221_pp0_iter5_reg <= data_31_V_read32_reg_4221_pp0_iter4_reg;
        data_31_V_read32_reg_4221_pp0_iter6_reg <= data_31_V_read32_reg_4221_pp0_iter5_reg;
        data_31_V_read32_reg_4221_pp0_iter7_reg <= data_31_V_read32_reg_4221_pp0_iter6_reg;
        data_31_V_read32_reg_4221_pp0_iter8_reg <= data_31_V_read32_reg_4221_pp0_iter7_reg;
        data_3_V_read_9_reg_5019 <= data_3_V_read_int_reg;
        data_3_V_read_9_reg_5019_pp0_iter1_reg <= data_3_V_read_9_reg_5019;
        data_3_V_read_9_reg_5019_pp0_iter2_reg <= data_3_V_read_9_reg_5019_pp0_iter1_reg;
        data_4_V_read_9_reg_4998 <= data_4_V_read_int_reg;
        data_4_V_read_9_reg_4998_pp0_iter1_reg <= data_4_V_read_9_reg_4998;
        data_4_V_read_9_reg_4998_pp0_iter2_reg <= data_4_V_read_9_reg_4998_pp0_iter1_reg;
        data_5_V_read_8_reg_4969 <= data_5_V_read_int_reg;
        data_5_V_read_8_reg_4969_pp0_iter1_reg <= data_5_V_read_8_reg_4969;
        data_5_V_read_8_reg_4969_pp0_iter2_reg <= data_5_V_read_8_reg_4969_pp0_iter1_reg;
        data_5_V_read_8_reg_4969_pp0_iter3_reg <= data_5_V_read_8_reg_4969_pp0_iter2_reg;
        data_6_V_read_8_reg_4944 <= data_6_V_read_int_reg;
        data_6_V_read_8_reg_4944_pp0_iter1_reg <= data_6_V_read_8_reg_4944;
        data_6_V_read_8_reg_4944_pp0_iter2_reg <= data_6_V_read_8_reg_4944_pp0_iter1_reg;
        data_6_V_read_8_reg_4944_pp0_iter3_reg <= data_6_V_read_8_reg_4944_pp0_iter2_reg;
        data_7_V_read_8_reg_4916 <= data_7_V_read_int_reg;
        data_7_V_read_8_reg_4916_pp0_iter1_reg <= data_7_V_read_8_reg_4916;
        data_7_V_read_8_reg_4916_pp0_iter2_reg <= data_7_V_read_8_reg_4916_pp0_iter1_reg;
        data_7_V_read_8_reg_4916_pp0_iter3_reg <= data_7_V_read_8_reg_4916_pp0_iter2_reg;
        data_8_V_read_7_reg_4887 <= data_8_V_read_int_reg;
        data_8_V_read_7_reg_4887_pp0_iter1_reg <= data_8_V_read_7_reg_4887;
        data_8_V_read_7_reg_4887_pp0_iter2_reg <= data_8_V_read_7_reg_4887_pp0_iter1_reg;
        data_8_V_read_7_reg_4887_pp0_iter3_reg <= data_8_V_read_7_reg_4887_pp0_iter2_reg;
        data_9_V_read_7_reg_4859 <= data_9_V_read_int_reg;
        data_9_V_read_7_reg_4859_pp0_iter1_reg <= data_9_V_read_7_reg_4859;
        data_9_V_read_7_reg_4859_pp0_iter2_reg <= data_9_V_read_7_reg_4859_pp0_iter1_reg;
        data_9_V_read_7_reg_4859_pp0_iter3_reg <= data_9_V_read_7_reg_4859_pp0_iter2_reg;
        data_9_V_read_7_reg_4859_pp0_iter4_reg <= data_9_V_read_7_reg_4859_pp0_iter3_reg;
        sub_ln703_105_reg_5226 <= sub_ln703_105_fu_489_p2;
        sub_ln703_113_reg_5247 <= sub_ln703_113_fu_533_p2;
        sub_ln703_114_reg_5253 <= sub_ln703_114_fu_549_p2;
        sub_ln703_117_reg_5259 <= sub_ln703_117_fu_554_p2;
        sub_ln703_126_reg_5274 <= sub_ln703_126_fu_574_p2;
        sub_ln703_129_reg_5279 <= sub_ln703_129_fu_579_p2;
        sub_ln703_133_reg_5284 <= sub_ln703_133_fu_584_p2;
        sub_ln703_138_reg_5325 <= sub_ln703_138_fu_816_p2;
        sub_ln703_141_reg_5330 <= sub_ln703_141_fu_835_p2;
        sub_ln703_143_reg_5335 <= sub_ln703_143_fu_844_p2;
        sub_ln703_144_reg_5340 <= sub_ln703_144_fu_858_p2;
        sub_ln703_145_reg_5345 <= sub_ln703_145_fu_863_p2;
        sub_ln703_149_reg_5350 <= sub_ln703_149_fu_901_p2;
        sub_ln703_154_reg_5355 <= sub_ln703_154_fu_920_p2;
        sub_ln703_161_reg_5365 <= sub_ln703_161_fu_960_p2;
        sub_ln703_162_reg_5370 <= sub_ln703_162_fu_980_p2;
        sub_ln703_166_reg_5375 <= sub_ln703_166_fu_1000_p2;
        sub_ln703_171_reg_5380 <= sub_ln703_171_fu_1015_p2;
        sub_ln703_173_reg_5385 <= sub_ln703_173_fu_1025_p2;
        sub_ln703_176_reg_5390 <= sub_ln703_176_fu_1040_p2;
        sub_ln703_180_reg_5395 <= sub_ln703_180_fu_1045_p2;
        sub_ln703_181_reg_5400 <= sub_ln703_181_fu_1050_p2;
        sub_ln703_182_reg_5410 <= sub_ln703_182_fu_1060_p2;
        sub_ln703_185_reg_5425 <= sub_ln703_185_fu_1095_p2;
        sub_ln703_187_reg_5440 <= sub_ln703_187_fu_1110_p2;
        sub_ln703_189_reg_5445 <= sub_ln703_189_fu_1115_p2;
        sub_ln703_191_reg_5450 <= sub_ln703_191_fu_1120_p2;
        sub_ln703_198_reg_5465 <= sub_ln703_198_fu_1146_p2;
        sub_ln703_199_reg_5470 <= sub_ln703_199_fu_1151_p2;
        sub_ln703_200_reg_5515 <= sub_ln703_200_fu_1326_p2;
        sub_ln703_203_reg_5520 <= sub_ln703_203_fu_1339_p2;
        sub_ln703_207_reg_5535 <= sub_ln703_207_fu_1384_p2;
        sub_ln703_212_reg_5540 <= sub_ln703_212_fu_1412_p2;
        sub_ln703_215_reg_5545 <= sub_ln703_215_fu_1441_p2;
        sub_ln703_229_reg_5560 <= sub_ln703_229_fu_1518_p2;
        sub_ln703_237_reg_5565 <= sub_ln703_237_fu_1571_p2;
        sub_ln703_238_reg_5570 <= sub_ln703_238_fu_1576_p2;
        sub_ln703_246_reg_5501 <= sub_ln703_246_fu_1193_p2;
        sub_ln703_252_reg_5575 <= sub_ln703_252_fu_1616_p2;
        sub_ln703_253_reg_5580 <= sub_ln703_253_fu_1621_p2;
        sub_ln703_254_reg_5585 <= sub_ln703_254_fu_1626_p2;
        sub_ln703_257_reg_5595 <= sub_ln703_257_fu_1641_p2;
        sub_ln703_261_reg_5600 <= sub_ln703_261_fu_1646_p2;
        sub_ln703_262_reg_5605 <= sub_ln703_262_fu_1651_p2;
        sub_ln703_263_reg_5610 <= sub_ln703_263_fu_1671_p2;
        sub_ln703_265_reg_5615 <= sub_ln703_265_fu_1676_p2;
        sub_ln703_266_reg_5620 <= sub_ln703_266_fu_1681_p2;
        sub_ln703_270_reg_5630 <= sub_ln703_270_fu_1695_p2;
        sub_ln703_272_reg_5635 <= sub_ln703_272_fu_1700_p2;
        sub_ln703_276_reg_5728 <= sub_ln703_276_fu_1918_p2;
        sub_ln703_278_reg_5650 <= sub_ln703_278_fu_1735_p2;
        sub_ln703_283_reg_5733 <= sub_ln703_283_fu_1975_p2;
        sub_ln703_288_reg_5738 <= sub_ln703_288_fu_2003_p2;
        sub_ln703_289_reg_5665 <= sub_ln703_289_fu_1750_p2;
        sub_ln703_290_reg_5670 <= sub_ln703_290_fu_1755_p2;
        sub_ln703_300_reg_5748 <= sub_ln703_300_fu_2075_p2;
        sub_ln703_302_reg_5758 <= sub_ln703_302_fu_2089_p2;
        sub_ln703_304_reg_5763 <= sub_ln703_304_fu_2099_p2;
        sub_ln703_309_reg_5773 <= sub_ln703_309_fu_2148_p2;
        sub_ln703_311_reg_5778 <= sub_ln703_311_fu_2173_p2;
        sub_ln703_318_reg_5783 <= sub_ln703_318_fu_2203_p2;
        sub_ln703_321_reg_5788 <= sub_ln703_321_fu_2218_p2;
        sub_ln703_323_reg_5798 <= sub_ln703_323_fu_2233_p2;
        sub_ln703_324_reg_5803 <= sub_ln703_324_fu_2238_p2;
        sub_ln703_325_reg_5808 <= sub_ln703_325_fu_2243_p2;
        sub_ln703_327_reg_5813 <= sub_ln703_327_fu_2248_p2;
        sub_ln703_328_reg_5818 <= sub_ln703_328_fu_2253_p2;
        sub_ln703_331_reg_5823 <= sub_ln703_331_fu_2258_p2;
        sub_ln703_332_reg_5828 <= sub_ln703_332_fu_2273_p2;
        sub_ln703_335_reg_5843 <= sub_ln703_335_fu_2302_p2;
        sub_ln703_343_reg_5853 <= sub_ln703_343_fu_2312_p2;
        sub_ln703_346_reg_5863 <= sub_ln703_346_fu_2332_p2;
        sub_ln703_356_reg_5921 <= sub_ln703_356_fu_2603_p2;
        sub_ln703_357_reg_5926 <= sub_ln703_357_fu_2608_p2;
        sub_ln703_361_reg_5936 <= sub_ln703_361_fu_2636_p2;
        sub_ln703_366_reg_5941 <= sub_ln703_366_fu_2684_p2;
        sub_ln703_369_reg_5946 <= sub_ln703_369_fu_2699_p2;
        sub_ln703_374_reg_5956 <= sub_ln703_374_fu_2728_p2;
        sub_ln703_375_reg_5966 <= sub_ln703_375_fu_2747_p2;
        sub_ln703_379_reg_5971 <= sub_ln703_379_fu_2781_p2;
        sub_ln703_381_reg_5976 <= sub_ln703_381_fu_2791_p2;
        sub_ln703_385_reg_5986 <= sub_ln703_385_fu_2811_p2;
        sub_ln703_386_reg_5991 <= sub_ln703_386_fu_2816_p2;
        sub_ln703_389_reg_5996 <= sub_ln703_389_fu_2839_p2;
        sub_ln703_392_reg_6001 <= sub_ln703_392_fu_2848_p2;
        sub_ln703_397_reg_6006 <= sub_ln703_397_fu_2863_p2;
        sub_ln703_402_reg_6016 <= sub_ln703_402_fu_2878_p2;
        sub_ln703_408_reg_6026 <= sub_ln703_408_fu_2893_p2;
        sub_ln703_409_reg_6031 <= sub_ln703_409_fu_2898_p2;
        sub_ln703_411_reg_6036 <= sub_ln703_411_fu_2903_p2;
        sub_ln703_416_reg_6046 <= sub_ln703_416_fu_2923_p2;
        sub_ln703_426_reg_6061 <= sub_ln703_426_fu_2938_p2;
        sub_ln703_428_reg_6108 <= sub_ln703_428_fu_3163_p2;
        sub_ln703_434_reg_6113 <= sub_ln703_434_fu_3199_p2;
        sub_ln703_448_reg_6118 <= sub_ln703_448_fu_3308_p2;
        sub_ln703_450_reg_6123 <= sub_ln703_450_fu_3318_p2;
        sub_ln703_451_reg_6143 <= sub_ln703_451_fu_3343_p2;
        sub_ln703_452_reg_6148 <= sub_ln703_452_fu_3348_p2;
        sub_ln703_453_reg_6153 <= sub_ln703_453_fu_3353_p2;
        sub_ln703_454_reg_6163 <= sub_ln703_454_fu_3368_p2;
        sub_ln703_455_reg_6168 <= sub_ln703_455_fu_3373_p2;
        sub_ln703_456_reg_6178 <= sub_ln703_456_fu_3388_p2;
        sub_ln703_457_reg_6183 <= sub_ln703_457_fu_3393_p2;
        sub_ln703_458_reg_6193 <= sub_ln703_458_fu_3408_p2;
        sub_ln703_459_reg_6198 <= sub_ln703_459_fu_3418_p2;
        sub_ln703_461_reg_6208 <= sub_ln703_461_fu_3438_p2;
        sub_ln703_469_reg_6218 <= sub_ln703_469_fu_3463_p2;
        sub_ln703_474_reg_6229 <= sub_ln703_474_fu_3482_p2;
        sub_ln703_486_reg_6244 <= sub_ln703_486_fu_3507_p2;
        sub_ln703_487_reg_6249 <= sub_ln703_487_fu_3512_p2;
        sub_ln703_491_reg_6254 <= sub_ln703_491_fu_3517_p2;
        sub_ln703_500_reg_6259 <= sub_ln703_500_fu_3522_p2;
        sub_ln703_73_reg_5059 <= sub_ln703_73_fu_286_p2;
        sub_ln703_74_reg_5065 <= sub_ln703_74_fu_292_p2;
        sub_ln703_74_reg_5065_pp0_iter2_reg <= sub_ln703_74_reg_5065;
        sub_ln703_76_reg_5071 <= sub_ln703_76_fu_300_p2;
        sub_ln703_76_reg_5071_pp0_iter2_reg <= sub_ln703_76_reg_5071;
        sub_ln703_77_reg_5084 <= sub_ln703_77_fu_308_p2;
        sub_ln703_79_reg_5125 <= sub_ln703_79_fu_337_p2;
        sub_ln703_89_reg_5166 <= sub_ln703_89_fu_402_p2;
        sub_ln703_91_reg_5172 <= sub_ln703_91_fu_411_p2;
        sub_ln703_93_reg_5200 <= sub_ln703_93_fu_442_p2;
        sub_ln703_94_reg_5205 <= sub_ln703_94_fu_446_p2;
        sub_ln703_96_reg_5210 <= sub_ln703_96_fu_456_p2;
        sub_ln703_reg_5046 <= sub_ln703_fu_274_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_511_fu_3847_p2;
        ap_return_10_int_reg <= acc_10_V_fu_3910_p2;
        ap_return_11_int_reg <= acc_11_V_fu_3915_p2;
        ap_return_12_int_reg <= acc_12_V_fu_3920_p2;
        ap_return_13_int_reg <= acc_13_V_fu_3925_p2;
        ap_return_14_int_reg <= acc_14_V_fu_3930_p2;
        ap_return_15_int_reg <= acc_15_V_fu_3935_p2;
        ap_return_16_int_reg <= acc_16_V_fu_3940_p2;
        ap_return_17_int_reg <= acc_17_V_fu_3953_p2;
        ap_return_18_int_reg <= acc_18_V_fu_3959_p2;
        ap_return_19_int_reg <= acc_19_V_fu_3964_p2;
        ap_return_1_int_reg <= acc_1_V_fu_3852_p2;
        ap_return_20_int_reg <= acc_20_V_fu_3969_p2;
        ap_return_21_int_reg <= acc_21_V_fu_3974_p2;
        ap_return_22_int_reg <= acc_22_V_fu_3979_p2;
        ap_return_23_int_reg <= acc_23_V_fu_3984_p2;
        ap_return_24_int_reg <= acc_24_V_fu_3989_p2;
        ap_return_25_int_reg <= acc_25_V_fu_3994_p2;
        ap_return_26_int_reg <= acc_26_V_fu_3999_p2;
        ap_return_27_int_reg <= acc_27_V_fu_4004_p2;
        ap_return_28_int_reg <= acc_28_V_fu_4009_p2;
        ap_return_29_int_reg <= acc_29_V_fu_4014_p2;
        ap_return_2_int_reg <= acc_2_V_fu_3857_p2;
        ap_return_30_int_reg <= acc_30_V_fu_4019_p2;
        ap_return_31_int_reg <= acc_31_V_fu_4024_p2;
        ap_return_3_int_reg <= acc_3_V_fu_3866_p2;
        ap_return_4_int_reg <= acc_4_V_fu_3879_p2;
        ap_return_5_int_reg <= acc_5_V_fu_3885_p2;
        ap_return_6_int_reg <= acc_6_V_fu_3890_p2;
        ap_return_7_int_reg <= acc_7_V_fu_3895_p2;
        ap_return_8_int_reg <= acc_8_V_fu_3900_p2;
        ap_return_9_int_reg <= acc_9_V_fu_3905_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_511_fu_3847_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_3852_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = acc_10_V_fu_3910_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = acc_11_V_fu_3915_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = acc_12_V_fu_3920_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = acc_13_V_fu_3925_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = acc_14_V_fu_3930_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = acc_15_V_fu_3935_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = acc_16_V_fu_3940_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = acc_17_V_fu_3953_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = acc_18_V_fu_3959_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = acc_19_V_fu_3964_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_3857_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = acc_20_V_fu_3969_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = acc_21_V_fu_3974_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = acc_22_V_fu_3979_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = acc_23_V_fu_3984_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = acc_24_V_fu_3989_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = acc_25_V_fu_3994_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = acc_26_V_fu_3999_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = acc_27_V_fu_4004_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = acc_28_V_fu_4009_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = acc_29_V_fu_4014_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_3866_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = acc_30_V_fu_4019_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = acc_31_V_fu_4024_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_3879_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = acc_5_V_fu_3885_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = acc_6_V_fu_3890_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = acc_7_V_fu_3895_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = acc_8_V_fu_3900_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = acc_9_V_fu_3905_p2;
    end
end

assign acc_10_V_fu_3910_p2 = (add_ln703_503_fu_3757_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_11_V_fu_3915_p2 = (sub_ln703_507_fu_3762_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_12_V_fu_3920_p2 = (sub_ln703_508_fu_3767_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_13_V_fu_3925_p2 = (sub_ln703_509_fu_3772_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_14_V_fu_3930_p2 = (add_ln703_504_fu_3777_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_15_V_fu_3935_p2 = (sub_ln703_510_fu_3781_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_16_V_fu_3940_p2 = (add_ln703_505_fu_3785_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_17_V_fu_3953_p2 = (add_ln703_527_fu_3949_p2 + add_ln703_526_fu_3945_p2);

assign acc_18_V_fu_3959_p2 = (sub_ln703_511_fu_3790_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_19_V_fu_3964_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_490_fu_3675_p2);

assign acc_1_V_fu_3852_p2 = (sub_ln703_501_fu_3728_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_20_V_fu_3969_p2 = (add_ln703_506_fu_3795_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_21_V_fu_3974_p2 = (add_ln703_507_fu_3799_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_22_V_fu_3979_p2 = (sub_ln703_512_fu_3804_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_23_V_fu_3984_p2 = (sub_ln703_513_fu_3809_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_24_V_fu_3989_p2 = (sub_ln703_514_fu_3814_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_25_V_fu_3994_p2 = (sub_ln703_515_fu_3819_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_26_V_fu_3999_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_497_fu_3704_p2);

assign acc_27_V_fu_4004_p2 = (sub_ln703_516_fu_3824_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_28_V_fu_4009_p2 = (sub_ln703_517_fu_3829_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_29_V_fu_4014_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_498_fu_3718_p2);

assign acc_2_V_fu_3857_p2 = (sub_ln703_502_fu_3732_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_30_V_fu_4019_p2 = (sub_ln703_518_fu_3834_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_31_V_fu_4024_p2 = (sub_ln703_519_fu_3839_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_3_V_fu_3866_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + add_ln703_514_fu_3862_p2);

assign acc_4_V_fu_3879_p2 = (add_ln703_518_fu_3875_p2 + add_ln703_517_fu_3871_p2);

assign acc_5_V_fu_3885_p2 = (sub_ln703_503_fu_3737_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_6_V_fu_3890_p2 = (sub_ln703_504_fu_3742_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_7_V_fu_3895_p2 = (sub_ln703_505_fu_3747_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_8_V_fu_3900_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_481_fu_3636_p2);

assign acc_9_V_fu_3905_p2 = (sub_ln703_506_fu_3752_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign add_ln703_200_fu_304_p2 = (add_ln703_reg_5052 + data_2_V_read_9_reg_5035);

assign add_ln703_201_fu_312_p2 = (sub_ln703_reg_5046 + data_2_V_read_9_reg_5035);

assign add_ln703_202_fu_316_p2 = (sub_ln703_73_reg_5059 + data_2_V_read_9_reg_5035);

assign add_ln703_203_fu_329_p2 = (sub_ln703_74_reg_5065 + data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign add_ln703_204_fu_320_p2 = (sub_ln703_75_fu_296_p2 + data_3_V_read_9_reg_5019);

assign add_ln703_205_fu_333_p2 = (add_ln703_200_reg_5077 + data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign add_ln703_206_fu_341_p2 = (sub_ln703_76_reg_5071 + data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign add_ln703_207_fu_325_p2 = (data_3_V_read_9_reg_5019 + data_4_V_read_9_reg_4998);

assign add_ln703_208_fu_345_p2 = (add_ln703_207_reg_5107 + sub_ln703_77_reg_5084);

assign add_ln703_209_fu_416_p2 = (add_ln703_205_reg_5119 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_210_fu_349_p2 = (add_ln703_204_reg_5101 + data_4_V_read_9_reg_4998_pp0_iter1_reg);

assign add_ln703_211_fu_420_p2 = (sub_ln703_82_fu_373_p2 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_212_fu_425_p2 = (add_ln703_203_reg_5113 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_213_fu_429_p2 = (add_ln703_207_reg_5107_pp0_iter2_reg + add_ln703_201_reg_5090_pp0_iter2_reg);

assign add_ln703_214_fu_433_p2 = (add_ln703_206_reg_5131 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_215_fu_605_p2 = (sub_ln703_89_reg_5166 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_216_fu_461_p2 = (sub_ln703_90_fu_406_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_217_fu_470_p2 = (add_ln703_210_reg_5143 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_218_fu_474_p2 = (add_ln703_211_fu_420_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_219_fu_479_p2 = (add_ln703_212_fu_425_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_220_fu_484_p2 = (sub_ln703_87_fu_393_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_221_fu_499_p2 = (add_ln703_208_reg_5137 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_222_fu_503_p2 = (data_5_V_read_8_reg_4969_pp0_iter2_reg + data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign add_ln703_223_fu_507_p2 = (add_ln703_222_fu_503_p2 + sub_ln703_85_fu_385_p2);

assign add_ln703_224_fu_645_p2 = (sub_ln703_96_reg_5210 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_225_fu_513_p2 = (sub_ln703_98_fu_466_p2 + data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign add_ln703_226_fu_518_p2 = (sub_ln703_79_reg_5125 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_227_fu_522_p2 = (add_ln703_222_fu_503_p2 + add_ln703_226_fu_518_p2);

assign add_ln703_228_fu_663_p2 = (sub_ln703_99_fu_613_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_229_fu_668_p2 = (sub_ln703_100_fu_617_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_230_fu_538_p2 = (sub_ln703_83_fu_377_p2 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_231_fu_543_p2 = (add_ln703_222_fu_503_p2 + add_ln703_230_fu_538_p2);

assign add_ln703_232_fu_673_p2 = (sub_ln703_101_fu_621_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_233_fu_353_p2 = (data_6_V_read_8_reg_4944_pp0_iter1_reg + data_7_V_read_8_reg_4916_pp0_iter1_reg);

assign add_ln703_234_fu_564_p2 = (add_ln703_233_reg_5149 + sub_ln703_95_fu_451_p2);

assign add_ln703_235_fu_701_p2 = (add_ln703_223_reg_5231 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_236_fu_710_p2 = (sub_ln703_111_fu_658_p2 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_237_fu_715_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + add_ln703_216_reg_5215);

assign add_ln703_238_fu_569_p2 = (add_ln703_233_reg_5149 + sub_ln703_94_fu_446_p2);

assign add_ln703_239_fu_750_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + sub_ln703_102_fu_625_p2);

assign add_ln703_240_fu_755_p2 = (sub_ln703_115_fu_678_p2 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_241_fu_765_p2 = (sub_ln703_117_reg_5259 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_242_fu_769_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + sub_ln703_107_fu_637_p2);

assign add_ln703_243_fu_774_p2 = (add_ln703_209_reg_5178 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_244_fu_778_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + add_ln703_243_fu_774_p2);

assign add_ln703_245_fu_783_p2 = (sub_ln703_114_reg_5253 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_246_fu_787_p2 = (sub_ln703_119_fu_687_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_247_fu_357_p2 = (data_7_V_read_8_reg_4916_pp0_iter1_reg + data_8_V_read_7_reg_4887_pp0_iter1_reg);

assign add_ln703_248_fu_801_p2 = (add_ln703_247_reg_5159_pp0_iter3_reg + sub_ln703_109_fu_649_p2);

assign add_ln703_249_fu_830_p2 = (sub_ln703_123_fu_719_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_250_fu_849_p2 = (sub_ln703_91_reg_5172 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_251_fu_589_p2 = (add_ln703_247_reg_5159 + data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign add_ln703_252_fu_853_p2 = (add_ln703_251_reg_5289 + add_ln703_250_fu_849_p2);

assign add_ln703_253_fu_873_p2 = (sub_ln703_105_reg_5226 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_254_fu_877_p2 = (add_ln703_247_reg_5159_pp0_iter3_reg + add_ln703_253_fu_873_p2);

assign add_ln703_255_fu_887_p2 = (add_ln703_214_reg_5194 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_256_fu_891_p2 = (add_ln703_251_reg_5289 + add_ln703_255_fu_887_p2);

assign add_ln703_257_fu_925_p2 = (sub_ln703_139_fu_821_p2 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_258_fu_593_p2 = (data_8_V_read_7_reg_4887_pp0_iter2_reg + data_9_V_read_7_reg_4859_pp0_iter2_reg);

assign add_ln703_259_fu_940_p2 = (add_ln703_258_reg_5295 + sub_ln703_124_fu_723_p2);

assign add_ln703_260_fu_950_p2 = (add_ln703_258_reg_5295 + sub_ln703_127_fu_732_p2);

assign add_ln703_261_fu_955_p2 = (add_ln703_258_reg_5295 + sub_ln703_131_fu_745_p2);

assign add_ln703_262_fu_965_p2 = (sub_ln703_104_fu_633_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_263_fu_970_p2 = (add_ln703_258_reg_5295 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_264_fu_974_p2 = (add_ln703_263_fu_970_p2 + add_ln703_262_fu_965_p2);

assign add_ln703_265_fu_1010_p2 = (sub_ln703_153_fu_915_p2 + data_10_V_read11_reg_4832_pp0_iter3_reg);

assign add_ln703_266_fu_1232_p2 = (sub_ln703_158_fu_1210_p2 + data_10_V_read11_reg_4832_pp0_iter4_reg);

assign add_ln703_267_fu_1055_p2 = (sub_ln703_164_fu_990_p2 + data_10_V_read11_reg_4832_pp0_iter3_reg);

assign add_ln703_268_fu_1065_p2 = (data_9_V_read_7_reg_4859_pp0_iter3_reg + data_10_V_read11_reg_4832_pp0_iter3_reg);

assign add_ln703_269_fu_1069_p2 = (add_ln703_268_fu_1065_p2 + sub_ln703_150_fu_906_p2);

assign add_ln703_270_fu_1255_p2 = (sub_ln703_169_fu_1222_p2 + data_11_V_read12_reg_4808_pp0_iter4_reg);

assign add_ln703_271_fu_1080_p2 = (sub_ln703_120_fu_691_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_272_fu_597_p2 = (data_10_V_read11_reg_4832_pp0_iter2_reg + data_11_V_read12_reg_4808_pp0_iter2_reg);

assign add_ln703_273_fu_1085_p2 = (add_ln703_272_reg_5304 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_274_fu_1089_p2 = (add_ln703_273_fu_1085_p2 + add_ln703_271_fu_1080_p2);

assign add_ln703_275_fu_1260_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + sub_ln703_154_reg_5355);

assign add_ln703_276_fu_1100_p2 = (sub_ln703_136_fu_806_p2 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_277_fu_1264_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + add_ln703_276_reg_5430);

assign add_ln703_278_fu_1105_p2 = (sub_ln703_137_fu_811_p2 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_279_fu_1268_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + add_ln703_278_reg_5435);

assign add_ln703_280_fu_1125_p2 = (sub_ln703_129_reg_5279 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_281_fu_1129_p2 = (add_ln703_273_fu_1085_p2 + add_ln703_280_fu_1125_p2);

assign add_ln703_282_fu_1135_p2 = (sub_ln703_130_fu_741_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_283_fu_1140_p2 = (add_ln703_273_fu_1085_p2 + add_ln703_282_fu_1135_p2);

assign add_ln703_284_fu_1296_p2 = (sub_ln703_145_reg_5345 + data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign add_ln703_285_fu_1300_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + add_ln703_284_fu_1296_p2);

assign add_ln703_286_fu_1305_p2 = (sub_ln703_180_reg_5395 + data_11_V_read12_reg_4808_pp0_iter4_reg);

assign add_ln703_287_fu_1354_p2 = (sub_ln703_186_fu_1272_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_288_fu_1156_p2 = (data_11_V_read12_reg_4808_pp0_iter3_reg + data_12_V_read13_reg_4778_pp0_iter3_reg);

assign add_ln703_289_fu_1359_p2 = (add_ln703_288_reg_5475 + sub_ln703_171_reg_5380);

assign add_ln703_290_fu_1367_p2 = (sub_ln703_189_reg_5445 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_291_fu_1371_p2 = (sub_ln703_190_fu_1281_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_292_fu_1376_p2 = (sub_ln703_191_reg_5450 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_293_fu_1380_p2 = (add_ln703_288_reg_5475 + sub_ln703_176_reg_5390);

assign add_ln703_294_fu_1397_p2 = (add_ln703_288_reg_5475 + sub_ln703_178_fu_1242_p2);

assign add_ln703_295_fu_1427_p2 = (sub_ln703_196_fu_1317_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_296_fu_1432_p2 = (sub_ln703_166_reg_5375 + data_10_V_read11_reg_4832_pp0_iter4_reg);

assign add_ln703_297_fu_1436_p2 = (add_ln703_288_reg_5475 + add_ln703_296_fu_1432_p2);

assign add_ln703_298_fu_1454_p2 = (sub_ln703_202_fu_1335_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_299_fu_1464_p2 = (sub_ln703_205_fu_1349_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_300_fu_1474_p2 = (sub_ln703_206_fu_1363_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_301_fu_1494_p2 = (sub_ln703_208_fu_1389_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_302_fu_1160_p2 = (sub_ln703_113_reg_5247 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_303_fu_1164_p2 = (add_ln703_258_reg_5295 + add_ln703_302_fu_1160_p2);

assign add_ln703_304_fu_601_p2 = (data_12_V_read13_reg_4778_pp0_iter2_reg + data_13_V_read14_reg_4745_pp0_iter2_reg);

assign add_ln703_305_fu_1169_p2 = (add_ln703_304_reg_5314 + add_ln703_272_reg_5304);

assign add_ln703_306_fu_1173_p2 = (add_ln703_305_fu_1169_p2 + add_ln703_303_fu_1164_p2);

assign add_ln703_307_fu_1504_p2 = (sub_ln703_210_fu_1402_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_308_fu_1509_p2 = (add_ln703_268_reg_5415 + sub_ln703_144_reg_5340);

assign add_ln703_309_fu_1179_p2 = (add_ln703_304_reg_5314 + data_11_V_read12_reg_4808_pp0_iter3_reg);

assign add_ln703_310_fu_1513_p2 = (add_ln703_309_reg_5484 + add_ln703_308_fu_1509_p2);

assign add_ln703_311_fu_1523_p2 = (sub_ln703_162_reg_5370 + data_10_V_read11_reg_4832_pp0_iter4_reg);

assign add_ln703_312_fu_1527_p2 = (add_ln703_309_reg_5484 + add_ln703_311_fu_1523_p2);

assign add_ln703_313_fu_1532_p2 = (sub_ln703_213_fu_1417_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_314_fu_1183_p2 = (data_13_V_read14_reg_4745_pp0_iter3_reg + data_14_V_read15_reg_4714_pp0_iter3_reg);

assign add_ln703_315_fu_1552_p2 = (add_ln703_314_reg_5490 + sub_ln703_201_fu_1331_p2);

assign add_ln703_316_fu_1187_p2 = (add_ln703_268_fu_1065_p2 + sub_ln703_135_fu_796_p2);

assign add_ln703_317_fu_1562_p2 = (add_ln703_314_reg_5490 + add_ln703_288_reg_5475);

assign add_ln703_318_fu_1566_p2 = (add_ln703_317_fu_1562_p2 + add_ln703_316_reg_5496);

assign add_ln703_319_fu_1591_p2 = (sub_ln703_223_fu_1479_p2 + data_14_V_read15_reg_4714_pp0_iter4_reg);

assign add_ln703_320_fu_1822_p2 = (sub_ln703_224_fu_1796_p2 + data_14_V_read15_reg_4714_pp0_iter5_reg);

assign add_ln703_321_fu_1636_p2 = (sub_ln703_236_fu_1557_p2 + data_15_V_read16_reg_4682_pp0_iter4_reg);

assign add_ln703_322_fu_1656_p2 = (sub_ln703_188_fu_1277_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_323_fu_1198_p2 = (data_14_V_read15_reg_4714_pp0_iter3_reg + data_15_V_read16_reg_4682_pp0_iter3_reg);

assign add_ln703_324_fu_1661_p2 = (add_ln703_323_reg_5506 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_325_fu_1665_p2 = (add_ln703_324_fu_1661_p2 + add_ln703_322_fu_1656_p2);

assign add_ln703_326_fu_1686_p2 = (add_ln703_323_reg_5506 + sub_ln703_228_fu_1499_p2);

assign add_ln703_327_fu_1887_p2 = (sub_ln703_250_fu_1844_p2 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_328_fu_1892_p2 = (sub_ln703_252_reg_5575 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_329_fu_1705_p2 = (sub_ln703_214_fu_1422_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_330_fu_1710_p2 = (add_ln703_323_reg_5506 + add_ln703_329_fu_1705_p2);

assign add_ln703_331_fu_1900_p2 = (sub_ln703_254_reg_5585 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_332_fu_1715_p2 = (sub_ln703_216_fu_1446_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_333_fu_1720_p2 = (add_ln703_323_reg_5506 + add_ln703_332_fu_1715_p2);

assign add_ln703_334_fu_1725_p2 = (add_ln703_323_reg_5506 + sub_ln703_234_fu_1547_p2);

assign add_ln703_335_fu_1730_p2 = (sub_ln703_256_fu_1631_p2 + data_16_V_read17_reg_4650_pp0_iter4_reg);

assign add_ln703_336_fu_1913_p2 = (sub_ln703_258_fu_1854_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_337_fu_1923_p2 = (sub_ln703_261_reg_5600 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_338_fu_1939_p2 = (sub_ln703_266_reg_5620 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_339_fu_1740_p2 = (sub_ln703_209_fu_1393_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_340_fu_1943_p2 = (data_15_V_read16_reg_4682_pp0_iter5_reg + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_341_fu_1947_p2 = (add_ln703_340_fu_1943_p2 + data_14_V_read15_reg_4714_pp0_iter5_reg);

assign add_ln703_342_fu_1952_p2 = (add_ln703_341_fu_1947_p2 + add_ln703_339_reg_5655);

assign add_ln703_343_fu_1745_p2 = (sub_ln703_268_fu_1691_p2 + data_16_V_read17_reg_4650_pp0_iter4_reg);

assign add_ln703_344_fu_1966_p2 = (sub_ln703_270_reg_5630 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_345_fu_1970_p2 = (sub_ln703_271_fu_1882_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_346_fu_1993_p2 = (sub_ln703_273_fu_1896_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_347_fu_1760_p2 = (data_16_V_read17_reg_4650_pp0_iter4_reg + data_17_V_read_8_reg_4621_pp0_iter4_reg);

assign add_ln703_348_fu_2017_p2 = (add_ln703_347_reg_5675 + sub_ln703_257_reg_5595);

assign add_ln703_349_fu_2021_p2 = (sub_ln703_219_fu_1788_p2 + data_14_V_read15_reg_4714_pp0_iter5_reg);

assign add_ln703_350_fu_2026_p2 = (add_ln703_347_reg_5675 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_351_fu_2030_p2 = (add_ln703_350_fu_2026_p2 + add_ln703_349_fu_2021_p2);

assign add_ln703_352_fu_2051_p2 = (sub_ln703_278_reg_5650 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_353_fu_2060_p2 = (add_ln703_347_reg_5675 + sub_ln703_264_fu_1867_p2);

assign add_ln703_354_fu_2080_p2 = (sub_ln703_281_fu_1957_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_355_fu_2114_p2 = (sub_ln703_290_reg_5670 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_356_fu_2118_p2 = (sub_ln703_235_fu_1812_p2 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_357_fu_1764_p2 = (data_17_V_read_8_reg_4621_pp0_iter4_reg + data_18_V_read_7_reg_4594_pp0_iter4_reg);

assign add_ln703_358_fu_2123_p2 = (add_ln703_357_reg_5683 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_359_fu_2127_p2 = (add_ln703_358_fu_2123_p2 + add_ln703_356_fu_2118_p2);

assign add_ln703_360_fu_2138_p2 = (sub_ln703_292_fu_2012_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_361_fu_2153_p2 = (sub_ln703_259_fu_1858_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_362_fu_2158_p2 = (add_ln703_357_reg_5683 + add_ln703_361_fu_2153_p2);

assign add_ln703_363_fu_2163_p2 = (sub_ln703_295_fu_2041_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_364_fu_2178_p2 = (sub_ln703_297_fu_2055_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_365_fu_2183_p2 = (sub_ln703_298_fu_2065_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_366_fu_2193_p2 = (sub_ln703_303_fu_2094_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_367_fu_2198_p2 = (sub_ln703_305_fu_2104_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_368_fu_2429_p2 = (add_ln703_357_reg_5683_pp0_iter6_reg + sub_ln703_288_reg_5738);

assign add_ln703_369_fu_2213_p2 = (sub_ln703_307_fu_2133_p2 + data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign add_ln703_370_fu_2437_p2 = (sub_ln703_309_reg_5773 + data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign add_ln703_371_fu_1768_p2 = (data_18_V_read_7_reg_4594_pp0_iter4_reg + data_19_V_read_7_reg_4567_pp0_iter4_reg);

assign add_ln703_372_fu_2228_p2 = (add_ln703_371_reg_5691 + sub_ln703_293_fu_2036_p2);

assign add_ln703_373_fu_2445_p2 = (sub_ln703_313_fu_2413_p2 + data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign add_ln703_374_fu_2263_p2 = (sub_ln703_284_fu_1980_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_375_fu_2268_p2 = (add_ln703_371_reg_5691 + add_ln703_374_fu_2263_p2);

assign add_ln703_376_fu_2278_p2 = (sub_ln703_287_fu_1998_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_377_fu_2283_p2 = (add_ln703_371_reg_5691 + add_ln703_376_fu_2278_p2);

assign add_ln703_378_fu_2288_p2 = (sub_ln703_289_reg_5665 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_379_fu_2292_p2 = (add_ln703_371_reg_5691 + add_ln703_378_fu_2288_p2);

assign add_ln703_380_fu_2297_p2 = (sub_ln703_319_fu_2208_p2 + data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign add_ln703_381_fu_2307_p2 = (sub_ln703_322_fu_2223_p2 + data_20_V_read21_reg_4539_pp0_iter5_reg);

assign add_ln703_382_fu_2486_p2 = (sub_ln703_325_reg_5808 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_383_fu_2490_p2 = (sub_ln703_326_fu_2441_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_384_fu_1772_p2 = (data_19_V_read_7_reg_4567_pp0_iter4_reg + data_20_V_read21_reg_4539_pp0_iter4_reg);

assign add_ln703_385_fu_2499_p2 = (add_ln703_384_reg_5701_pp0_iter6_reg + sub_ln703_312_fu_2409_p2);

assign add_ln703_386_fu_2514_p2 = (sub_ln703_331_reg_5823 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_387_fu_2518_p2 = (add_ln703_384_reg_5701_pp0_iter6_reg + sub_ln703_317_fu_2425_p2);

assign add_ln703_388_fu_2317_p2 = (sub_ln703_285_fu_1984_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_389_fu_2322_p2 = (add_ln703_384_reg_5701 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_390_fu_2326_p2 = (add_ln703_389_fu_2322_p2 + add_ln703_388_fu_2317_p2);

assign add_ln703_391_fu_2527_p2 = (sub_ln703_334_fu_2464_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_392_fu_2540_p2 = (sub_ln703_336_fu_2469_p2 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_393_fu_2559_p2 = (sub_ln703_294_fu_2405_p2 + data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign add_ln703_394_fu_1776_p2 = (data_20_V_read21_reg_4539_pp0_iter4_reg + data_21_V_read22_reg_4512_pp0_iter4_reg);

assign add_ln703_395_fu_2564_p2 = (add_ln703_394_reg_5710_pp0_iter6_reg + data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign add_ln703_396_fu_2568_p2 = (add_ln703_395_fu_2564_p2 + add_ln703_393_fu_2559_p2);

assign add_ln703_397_fu_2599_p2 = (add_ln703_394_reg_5710_pp0_iter6_reg + sub_ln703_328_reg_5818);

assign add_ln703_398_fu_2337_p2 = (add_ln703_347_reg_5675 + sub_ln703_267_fu_1872_p2);

assign add_ln703_399_fu_2342_p2 = (add_ln703_394_reg_5710 + add_ln703_371_reg_5691);

assign add_ln703_400_fu_2346_p2 = (add_ln703_399_fu_2342_p2 + add_ln703_398_fu_2337_p2);

assign add_ln703_401_fu_2623_p2 = (sub_ln703_343_reg_5853 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_402_fu_2631_p2 = (sub_ln703_344_fu_2523_p2 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_403_fu_2645_p2 = (sub_ln703_320_fu_2433_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_404_fu_1780_p2 = (data_21_V_read22_reg_4512_pp0_iter4_reg + data_22_V_read23_reg_4483_pp0_iter4_reg);

assign add_ln703_405_fu_2650_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_403_fu_2645_p2);

assign add_ln703_406_fu_2655_p2 = (sub_ln703_347_fu_2536_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_407_fu_2675_p2 = (sub_ln703_323_reg_5798 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_408_fu_2679_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_407_fu_2675_p2);

assign add_ln703_409_fu_2704_p2 = (sub_ln703_354_fu_2589_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_410_fu_2709_p2 = (sub_ln703_355_fu_2594_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_411_fu_2352_p2 = (add_ln703_371_reg_5691 + sub_ln703_299_fu_2070_p2);

assign add_ln703_412_fu_2357_p2 = (add_ln703_404_reg_5718 + data_20_V_read21_reg_4539_pp0_iter5_reg);

assign add_ln703_413_fu_2361_p2 = (add_ln703_412_fu_2357_p2 + add_ln703_411_fu_2352_p2);

assign add_ln703_414_fu_2367_p2 = (sub_ln703_315_fu_2188_p2 + data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign add_ln703_415_fu_2372_p2 = (add_ln703_412_fu_2357_p2 + add_ln703_414_fu_2367_p2);

assign add_ln703_416_fu_2733_p2 = (add_ln703_357_reg_5683_pp0_iter6_reg + sub_ln703_283_reg_5733);

assign add_ln703_417_fu_2737_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_384_reg_5701_pp0_iter6_reg);

assign add_ln703_418_fu_2741_p2 = (add_ln703_417_fu_2737_p2 + add_ln703_416_fu_2733_p2);

assign add_ln703_419_fu_2757_p2 = (sub_ln703_332_reg_5828 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_420_fu_2761_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_419_fu_2757_p2);

assign add_ln703_421_fu_2766_p2 = (sub_ln703_333_fu_2460_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_422_fu_2771_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_421_fu_2766_p2);

assign add_ln703_423_fu_2993_p2 = (sub_ln703_361_reg_5936 + data_22_V_read23_reg_4483_pp0_iter7_reg);

assign add_ln703_424_fu_2806_p2 = (sub_ln703_367_fu_2689_p2 + data_23_V_read24_reg_4451_pp0_iter6_reg);

assign add_ln703_425_fu_3001_p2 = (sub_ln703_369_reg_5946 + data_23_V_read24_reg_4451_pp0_iter7_reg);

assign add_ln703_426_fu_2378_p2 = (sub_ln703_244_fu_1827_p2 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_427_fu_2383_p2 = (add_ln703_358_fu_2123_p2 + add_ln703_426_fu_2378_p2);

assign add_ln703_428_fu_2389_p2 = (data_22_V_read23_reg_4483_pp0_iter5_reg + data_23_V_read24_reg_4451_pp0_iter5_reg);

assign add_ln703_429_fu_2825_p2 = (add_ln703_428_reg_5888 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_430_fu_2829_p2 = (add_ln703_429_fu_2825_p2 + add_ln703_384_reg_5701_pp0_iter6_reg);

assign add_ln703_431_fu_2834_p2 = (add_ln703_430_fu_2829_p2 + add_ln703_427_reg_5883);

assign add_ln703_432_fu_3014_p2 = (sub_ln703_374_reg_5956 + data_23_V_read24_reg_4451_pp0_iter7_reg);

assign add_ln703_433_fu_3036_p2 = (sub_ln703_379_reg_5971 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_434_fu_2873_p2 = (sub_ln703_380_fu_2786_p2 + data_24_V_read25_reg_4421_pp0_iter6_reg);

assign add_ln703_435_fu_2393_p2 = (data_23_V_read24_reg_4451_pp0_iter5_reg + data_24_V_read25_reg_4421_pp0_iter5_reg);

assign add_ln703_436_fu_2883_p2 = (add_ln703_435_reg_5894 + sub_ln703_365_fu_2670_p2);

assign add_ln703_437_fu_3053_p2 = (sub_ln703_385_reg_5986 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_438_fu_2888_p2 = (add_ln703_435_reg_5894 + sub_ln703_370_fu_2714_p2);

assign add_ln703_439_fu_3075_p2 = (sub_ln703_390_fu_3009_p2 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_440_fu_2908_p2 = (add_ln703_394_reg_5710_pp0_iter6_reg + sub_ln703_330_fu_2455_p2);

assign add_ln703_441_fu_2913_p2 = (add_ln703_435_reg_5894 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_442_fu_2917_p2 = (add_ln703_441_fu_2913_p2 + add_ln703_440_fu_2908_p2);

assign add_ln703_443_fu_3099_p2 = (sub_ln703_397_reg_6006 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_444_fu_2928_p2 = (sub_ln703_400_fu_2868_p2 + data_24_V_read25_reg_4421_pp0_iter6_reg);

assign add_ln703_445_fu_3122_p2 = (sub_ln703_402_reg_6016 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_446_fu_2397_p2 = (data_24_V_read25_reg_4421_pp0_iter5_reg + data_25_V_read26_reg_4391_pp0_iter5_reg);

assign add_ln703_447_fu_2933_p2 = (add_ln703_446_reg_5901 + sub_ln703_383_fu_2801_p2);

assign add_ln703_448_fu_3150_p2 = (sub_ln703_408_reg_6026 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_449_fu_3158_p2 = (sub_ln703_410_fu_3071_p2 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_450_fu_3168_p2 = (sub_ln703_357_reg_5926 + data_22_V_read23_reg_4483_pp0_iter7_reg);

assign add_ln703_451_fu_2943_p2 = (add_ln703_446_reg_5901 + data_23_V_read24_reg_4451_pp0_iter6_reg);

assign add_ln703_452_fu_3172_p2 = (add_ln703_451_reg_6066 + add_ln703_450_fu_3168_p2);

assign add_ln703_453_fu_3218_p2 = (sub_ln703_420_fu_3117_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_454_fu_3232_p2 = (sub_ln703_424_fu_3140_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_455_fu_3237_p2 = (data_25_V_read26_reg_4391_pp0_iter7_reg + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_456_fu_3241_p2 = (add_ln703_455_fu_3237_p2 + sub_ln703_405_fu_3057_p2);

assign add_ln703_457_fu_3281_p2 = (sub_ln703_431_fu_3185_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_458_fu_3286_p2 = (add_ln703_455_fu_3237_p2 + sub_ln703_413_fu_3084_p2);

assign add_ln703_459_fu_3292_p2 = (add_ln703_455_fu_3237_p2 + sub_ln703_415_fu_3094_p2);

assign add_ln703_460_fu_3303_p2 = (sub_ln703_433_fu_3194_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_461_fu_3323_p2 = (sub_ln703_438_fu_3223_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_462_fu_2401_p2 = (data_26_V_read27_reg_4365_pp0_iter5_reg + data_27_V_read_8_reg_4342_pp0_iter5_reg);

assign add_ln703_463_fu_3328_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + sub_ln703_421_fu_3126_p2);

assign add_ln703_464_fu_3333_p2 = (sub_ln703_439_fu_3228_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_465_fu_3338_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + sub_ln703_422_fu_3130_p2);

assign add_ln703_466_fu_3358_p2 = (sub_ln703_407_fu_3066_p2 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_467_fu_3363_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + add_ln703_466_fu_3358_p2);

assign add_ln703_468_fu_3378_p2 = (sub_ln703_445_fu_3271_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_469_fu_3383_p2 = (sub_ln703_446_fu_3276_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_470_fu_3398_p2 = (sub_ln703_414_fu_3089_p2 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_471_fu_3403_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + add_ln703_470_fu_3398_p2);

assign add_ln703_472_fu_3413_p2 = (sub_ln703_447_fu_3298_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_473_fu_3423_p2 = (sub_ln703_398_fu_3026_p2 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_474_fu_3428_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_475_fu_3432_p2 = (add_ln703_474_fu_3428_p2 + add_ln703_473_fu_3423_p2);

assign add_ln703_476_fu_3531_p2 = (add_ln703_462_reg_5909_pp0_iter8_reg + sub_ln703_434_reg_6113);

assign add_ln703_477_fu_2947_p2 = (sub_ln703_345_fu_2532_p2 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_478_fu_2952_p2 = (add_ln703_428_reg_5888 + add_ln703_477_fu_2947_p2);

assign add_ln703_479_fu_2957_p2 = (add_ln703_462_reg_5909 + add_ln703_446_reg_5901);

assign add_ln703_480_fu_2961_p2 = (add_ln703_479_fu_2957_p2 + add_ln703_478_fu_2952_p2);

assign add_ln703_481_fu_3443_p2 = (sub_ln703_423_fu_3135_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_482_fu_2967_p2 = (data_27_V_read_8_reg_4342_pp0_iter6_reg + data_28_V_read_7_reg_4313_pp0_iter6_reg);

assign add_ln703_483_fu_3448_p2 = (add_ln703_482_reg_6077 + add_ln703_481_fu_3443_p2);

assign add_ln703_484_fu_3555_p2 = (sub_ln703_452_reg_6148 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_485_fu_3559_p2 = (sub_ln703_453_reg_6153 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_486_fu_3453_p2 = (add_ln703_482_reg_6077 + sub_ln703_442_fu_3256_p2);

assign add_ln703_487_fu_3458_p2 = (add_ln703_482_reg_6077 + sub_ln703_443_fu_3261_p2);

assign add_ln703_488_fu_3571_p2 = (sub_ln703_455_reg_6168 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_489_fu_3468_p2 = (sub_ln703_430_fu_3181_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_490_fu_3473_p2 = (add_ln703_482_reg_6077 + add_ln703_489_fu_3468_p2);

assign add_ln703_491_fu_2971_p2 = (add_ln703_446_reg_5901 + sub_ln703_395_fu_2853_p2);

assign add_ln703_492_fu_3478_p2 = (add_ln703_482_reg_6077 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_493_fu_3595_p2 = (add_ln703_492_reg_6223 + add_ln703_491_reg_6087_pp0_iter8_reg);

assign add_ln703_494_fu_3487_p2 = (sub_ln703_435_fu_3204_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_495_fu_3492_p2 = (add_ln703_482_reg_6077 + add_ln703_494_fu_3487_p2);

assign add_ln703_496_fu_3497_p2 = (data_28_V_read_7_reg_4313_pp0_iter7_reg + data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign add_ln703_497_fu_3501_p2 = (add_ln703_496_fu_3497_p2 + sub_ln703_449_fu_3313_p2);

assign add_ln703_498_fu_3616_p2 = (sub_ln703_460_fu_3535_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_499_fu_3631_p2 = (sub_ln703_464_fu_3547_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_500_fu_3655_p2 = (sub_ln703_466_fu_3563_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_501_fu_3708_p2 = (sub_ln703_475_fu_3599_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_502_fu_3713_p2 = (sub_ln703_476_fu_3603_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_503_fu_3757_p2 = (sub_ln703_483_fu_3645_p2 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_504_fu_3777_p2 = (sub_ln703_486_reg_6244 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_505_fu_3785_p2 = (sub_ln703_488_fu_3665_p2 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_506_fu_3795_p2 = (sub_ln703_491_reg_6254 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_507_fu_3799_p2 = (sub_ln703_492_fu_3679_p2 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_508_fu_3843_p2 = (sub_ln703_448_reg_6118 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_509_fu_2976_p2 = (data_30_V_read31_reg_4250_pp0_iter6_reg + data_31_V_read32_reg_4221_pp0_iter6_reg);

assign add_ln703_510_fu_3527_p2 = (add_ln703_509_reg_6092 + data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign add_ln703_511_fu_3847_p2 = (add_ln703_510_reg_6264 + add_ln703_508_fu_3843_p2);

assign add_ln703_514_fu_3862_p2 = (sub_ln703_461_reg_6208 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_516_fu_2980_p2 = (sub_ln703_349_fu_2549_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_517_fu_3871_p2 = (add_ln703_451_reg_6066_pp0_iter8_reg + add_ln703_516_reg_6103_pp0_iter8_reg);

assign add_ln703_518_fu_3875_p2 = (add_ln703_510_reg_6264 + add_ln703_492_reg_6223);

assign add_ln703_526_fu_3945_p2 = (add_ln703_462_reg_5909_pp0_iter8_reg + sub_ln703_428_reg_6108);

assign add_ln703_527_fu_3949_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + add_ln703_496_reg_6234);

assign add_ln703_fu_280_p2 = (data_0_V_read_int_reg + data_1_V_read_int_reg);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign sub_ln703_100_fu_617_p2 = (add_ln703_210_reg_5143_pp0_iter3_reg - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_101_fu_621_p2 = (add_ln703_213_reg_5189 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_102_fu_625_p2 = (sub_ln703_89_reg_5166 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_103_fu_629_p2 = (add_ln703_214_reg_5194 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_104_fu_633_p2 = (add_ln703_211_reg_5184 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_105_fu_489_p2 = (sub_ln703_92_fu_437_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_106_fu_494_p2 = (add_ln703_212_fu_425_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_107_fu_637_p2 = (sub_ln703_93_reg_5200 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_108_fu_641_p2 = (sub_ln703_94_reg_5205 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_109_fu_649_p2 = (add_ln703_215_fu_605_p2 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_110_fu_654_p2 = (add_ln703_216_reg_5215 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_111_fu_658_p2 = (sub_ln703_97_fu_609_p2 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_112_fu_528_p2 = (add_ln703_217_fu_470_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_113_fu_533_p2 = (add_ln703_218_fu_474_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_114_fu_549_p2 = (add_ln703_219_fu_479_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_115_fu_678_p2 = (sub_ln703_103_fu_629_p2 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_116_fu_683_p2 = (add_ln703_220_reg_5221 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_117_fu_554_p2 = (sub_ln703_106_fu_494_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_118_fu_559_p2 = (add_ln703_221_fu_499_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_119_fu_687_p2 = (add_ln703_223_reg_5231 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_120_fu_691_p2 = (sub_ln703_108_fu_641_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_121_fu_696_p2 = (add_ln703_224_fu_645_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_122_fu_705_p2 = (sub_ln703_110_fu_654_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_123_fu_719_p2 = (add_ln703_225_reg_5237 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_124_fu_723_p2 = (add_ln703_227_reg_5242 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_125_fu_727_p2 = (add_ln703_228_fu_663_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_126_fu_574_p2 = (sub_ln703_112_fu_528_p2 - data_7_V_read_8_reg_4916_pp0_iter2_reg);

assign sub_ln703_127_fu_732_p2 = (sub_ln703_113_reg_5247 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_128_fu_736_p2 = (add_ln703_229_fu_668_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_129_fu_579_p2 = (add_ln703_231_fu_543_p2 - data_7_V_read_8_reg_4916_pp0_iter2_reg);

assign sub_ln703_130_fu_741_p2 = (sub_ln703_114_reg_5253 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_131_fu_745_p2 = (add_ln703_232_fu_673_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_132_fu_760_p2 = (sub_ln703_116_fu_683_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_133_fu_584_p2 = (sub_ln703_118_fu_559_p2 - data_7_V_read_8_reg_4916_pp0_iter2_reg);

assign sub_ln703_134_fu_792_p2 = (add_ln703_234_reg_5264 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_135_fu_796_p2 = (sub_ln703_121_fu_696_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_136_fu_806_p2 = (add_ln703_235_fu_701_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_137_fu_811_p2 = (sub_ln703_122_fu_705_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_138_fu_816_p2 = (add_ln703_236_fu_710_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_139_fu_821_p2 = (add_ln703_237_fu_715_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_140_fu_826_p2 = (add_ln703_238_reg_5269 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_141_fu_835_p2 = (sub_ln703_125_fu_727_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_142_fu_840_p2 = (sub_ln703_126_reg_5274 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_143_fu_844_p2 = (sub_ln703_128_fu_736_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_144_fu_858_p2 = (add_ln703_239_fu_750_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_145_fu_863_p2 = (add_ln703_240_fu_755_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_146_fu_868_p2 = (sub_ln703_132_fu_760_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_147_fu_882_p2 = (add_ln703_241_fu_765_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_148_fu_896_p2 = (add_ln703_242_fu_769_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_149_fu_901_p2 = (add_ln703_244_fu_778_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_150_fu_906_p2 = (add_ln703_245_fu_783_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_151_fu_911_p2 = (sub_ln703_133_reg_5284 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_152_fu_1202_p2 = (add_ln703_246_reg_5320 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_153_fu_915_p2 = (sub_ln703_134_fu_792_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_154_fu_920_p2 = (add_ln703_248_fu_801_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_155_fu_1206_p2 = (sub_ln703_138_reg_5325 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_156_fu_930_p2 = (sub_ln703_140_fu_826_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_157_fu_935_p2 = (add_ln703_249_fu_830_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_158_fu_1210_p2 = (sub_ln703_141_reg_5330 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_159_fu_945_p2 = (sub_ln703_142_fu_840_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_160_fu_1214_p2 = (sub_ln703_143_reg_5335 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_161_fu_960_p2 = (add_ln703_252_fu_853_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_162_fu_980_p2 = (sub_ln703_146_fu_868_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_163_fu_985_p2 = (add_ln703_254_fu_877_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_164_fu_990_p2 = (sub_ln703_147_fu_882_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_165_fu_995_p2 = (add_ln703_256_fu_891_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_166_fu_1000_p2 = (sub_ln703_148_fu_896_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_167_fu_1218_p2 = (sub_ln703_149_reg_5350 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_168_fu_1005_p2 = (sub_ln703_151_fu_911_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_169_fu_1222_p2 = (sub_ln703_152_fu_1202_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_170_fu_1227_p2 = (sub_ln703_155_fu_1206_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_171_fu_1015_p2 = (add_ln703_257_fu_925_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_172_fu_1020_p2 = (sub_ln703_156_fu_930_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_173_fu_1025_p2 = (sub_ln703_157_fu_935_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_174_fu_1030_p2 = (add_ln703_259_fu_940_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_175_fu_1035_p2 = (sub_ln703_159_fu_945_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_176_fu_1040_p2 = (add_ln703_260_fu_950_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_177_fu_1237_p2 = (sub_ln703_160_fu_1214_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_178_fu_1242_p2 = (add_ln703_261_reg_5360 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_179_fu_1246_p2 = (sub_ln703_161_reg_5365 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_180_fu_1045_p2 = (add_ln703_264_fu_974_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_181_fu_1050_p2 = (sub_ln703_163_fu_985_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_182_fu_1060_p2 = (sub_ln703_165_fu_995_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_183_fu_1250_p2 = (sub_ln703_167_fu_1218_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_184_fu_1075_p2 = (sub_ln703_168_fu_1005_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_185_fu_1095_p2 = (add_ln703_265_fu_1010_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_186_fu_1272_p2 = (sub_ln703_170_fu_1227_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_187_fu_1110_p2 = (sub_ln703_172_fu_1020_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_188_fu_1277_p2 = (sub_ln703_173_reg_5385 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_189_fu_1115_p2 = (sub_ln703_174_fu_1030_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_190_fu_1281_p2 = (add_ln703_266_fu_1232_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_191_fu_1120_p2 = (sub_ln703_175_fu_1035_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_192_fu_1286_p2 = (sub_ln703_177_fu_1237_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_193_fu_1291_p2 = (sub_ln703_179_fu_1246_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_194_fu_1309_p2 = (sub_ln703_181_reg_5400 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_195_fu_1313_p2 = (add_ln703_267_reg_5405 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_196_fu_1317_p2 = (sub_ln703_182_reg_5410 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_197_fu_1321_p2 = (sub_ln703_183_fu_1250_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_198_fu_1146_p2 = (add_ln703_269_fu_1069_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_199_fu_1151_p2 = (sub_ln703_184_fu_1075_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_200_fu_1326_p2 = (add_ln703_270_fu_1255_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_201_fu_1331_p2 = (add_ln703_274_reg_5420 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_202_fu_1335_p2 = (sub_ln703_185_reg_5425 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_203_fu_1339_p2 = (add_ln703_275_fu_1260_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_204_fu_1344_p2 = (add_ln703_277_fu_1264_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_205_fu_1349_p2 = (add_ln703_279_fu_1268_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_206_fu_1363_p2 = (sub_ln703_187_reg_5440 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_207_fu_1384_p2 = (sub_ln703_192_fu_1286_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_208_fu_1389_p2 = (add_ln703_281_reg_5455 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_209_fu_1393_p2 = (add_ln703_283_reg_5460 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_210_fu_1402_p2 = (sub_ln703_193_fu_1291_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_211_fu_1407_p2 = (add_ln703_285_fu_1300_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_212_fu_1412_p2 = (add_ln703_286_fu_1305_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_213_fu_1417_p2 = (sub_ln703_194_fu_1309_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_214_fu_1422_p2 = (sub_ln703_195_fu_1313_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_215_fu_1441_p2 = (sub_ln703_197_fu_1321_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_216_fu_1446_p2 = (sub_ln703_198_reg_5465 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_217_fu_1450_p2 = (sub_ln703_199_reg_5470 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_218_fu_1784_p2 = (sub_ln703_200_reg_5515 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_219_fu_1788_p2 = (sub_ln703_203_reg_5520 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_220_fu_1459_p2 = (sub_ln703_204_fu_1344_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_221_fu_1792_p2 = (add_ln703_287_reg_5525 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_222_fu_1469_p2 = (add_ln703_289_fu_1359_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_223_fu_1479_p2 = (add_ln703_290_fu_1367_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_224_fu_1796_p2 = (add_ln703_291_reg_5530 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_225_fu_1484_p2 = (add_ln703_292_fu_1376_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_226_fu_1489_p2 = (add_ln703_293_fu_1380_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_227_fu_1800_p2 = (sub_ln703_207_reg_5535 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_228_fu_1499_p2 = (add_ln703_294_fu_1397_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_229_fu_1518_p2 = (sub_ln703_211_fu_1407_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_230_fu_1804_p2 = (sub_ln703_212_reg_5540 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_231_fu_1537_p2 = (add_ln703_295_fu_1427_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_232_fu_1542_p2 = (add_ln703_297_fu_1436_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_233_fu_1808_p2 = (sub_ln703_215_reg_5545 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_234_fu_1547_p2 = (sub_ln703_217_fu_1450_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_235_fu_1812_p2 = (sub_ln703_218_fu_1784_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_236_fu_1557_p2 = (add_ln703_298_fu_1454_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_237_fu_1571_p2 = (sub_ln703_220_fu_1459_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_238_fu_1576_p2 = (add_ln703_299_fu_1464_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_239_fu_1817_p2 = (sub_ln703_221_fu_1792_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_240_fu_1581_p2 = (sub_ln703_222_fu_1469_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_241_fu_1586_p2 = (add_ln703_300_fu_1474_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_242_fu_1596_p2 = (sub_ln703_225_fu_1484_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_243_fu_1601_p2 = (sub_ln703_226_fu_1489_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_244_fu_1827_p2 = (sub_ln703_227_fu_1800_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_245_fu_1832_p2 = (add_ln703_301_reg_5550 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_246_fu_1193_p2 = (add_ln703_306_fu_1173_p2 - data_14_V_read15_reg_4714_pp0_iter3_reg);

assign sub_ln703_247_fu_1836_p2 = (add_ln703_307_reg_5555 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_248_fu_1606_p2 = (add_ln703_310_fu_1513_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_249_fu_1840_p2 = (sub_ln703_229_reg_5560 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_250_fu_1844_p2 = (sub_ln703_230_fu_1804_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_251_fu_1611_p2 = (add_ln703_312_fu_1527_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_252_fu_1616_p2 = (add_ln703_313_fu_1532_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_253_fu_1621_p2 = (sub_ln703_231_fu_1537_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_254_fu_1626_p2 = (sub_ln703_232_fu_1542_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_255_fu_1849_p2 = (sub_ln703_233_fu_1808_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_256_fu_1631_p2 = (add_ln703_315_fu_1552_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_257_fu_1641_p2 = (add_ln703_318_fu_1566_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_258_fu_1854_p2 = (sub_ln703_237_reg_5565 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_259_fu_1858_p2 = (sub_ln703_238_reg_5570 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_260_fu_1862_p2 = (sub_ln703_239_fu_1817_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_261_fu_1646_p2 = (sub_ln703_240_fu_1581_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_262_fu_1651_p2 = (sub_ln703_241_fu_1586_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_263_fu_1671_p2 = (add_ln703_319_fu_1591_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_264_fu_1867_p2 = (add_ln703_320_fu_1822_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_265_fu_1676_p2 = (sub_ln703_242_fu_1596_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_266_fu_1681_p2 = (sub_ln703_243_fu_1601_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_267_fu_1872_p2 = (sub_ln703_245_fu_1832_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_268_fu_1691_p2 = (sub_ln703_246_reg_5501 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_269_fu_1877_p2 = (sub_ln703_247_fu_1836_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_270_fu_1695_p2 = (sub_ln703_248_fu_1606_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_271_fu_1882_p2 = (sub_ln703_249_fu_1840_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_272_fu_1700_p2 = (sub_ln703_251_fu_1611_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_273_fu_1896_p2 = (sub_ln703_253_reg_5580 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_274_fu_1904_p2 = (sub_ln703_255_fu_1849_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_275_fu_1909_p2 = (add_ln703_321_reg_5590 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_276_fu_1918_p2 = (sub_ln703_260_fu_1862_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_277_fu_1927_p2 = (sub_ln703_262_reg_5605 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_278_fu_1735_p2 = (add_ln703_325_fu_1665_p2 - data_16_V_read17_reg_4650_pp0_iter4_reg);

assign sub_ln703_279_fu_1931_p2 = (sub_ln703_263_reg_5610 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_280_fu_1935_p2 = (sub_ln703_265_reg_5615 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_281_fu_1957_p2 = (add_ln703_326_reg_5625 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_282_fu_1961_p2 = (sub_ln703_269_fu_1877_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_283_fu_1975_p2 = (add_ln703_327_fu_1887_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_284_fu_1980_p2 = (sub_ln703_272_reg_5635 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_285_fu_1984_p2 = (add_ln703_328_fu_1892_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_286_fu_1989_p2 = (add_ln703_330_reg_5640 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_287_fu_1998_p2 = (add_ln703_331_fu_1900_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_288_fu_2003_p2 = (sub_ln703_274_fu_1904_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_289_fu_1750_p2 = (add_ln703_333_fu_1720_p2 - data_16_V_read17_reg_4650_pp0_iter4_reg);

assign sub_ln703_290_fu_1755_p2 = (add_ln703_334_fu_1725_p2 - data_16_V_read17_reg_4650_pp0_iter4_reg);

assign sub_ln703_291_fu_2008_p2 = (add_ln703_335_reg_5645 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_292_fu_2012_p2 = (sub_ln703_275_fu_1909_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_293_fu_2036_p2 = (add_ln703_336_fu_1913_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_294_fu_2405_p2 = (sub_ln703_276_reg_5728 - data_17_V_read_8_reg_4621_pp0_iter6_reg);

assign sub_ln703_295_fu_2041_p2 = (add_ln703_337_fu_1923_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_296_fu_2046_p2 = (sub_ln703_277_fu_1927_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_297_fu_2055_p2 = (sub_ln703_279_fu_1931_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_298_fu_2065_p2 = (sub_ln703_280_fu_1935_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_299_fu_2070_p2 = (add_ln703_338_fu_1939_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_300_fu_2075_p2 = (add_ln703_342_fu_1952_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_301_fu_2085_p2 = (add_ln703_343_reg_5660 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_302_fu_2089_p2 = (sub_ln703_282_fu_1961_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_303_fu_2094_p2 = (add_ln703_344_fu_1966_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_304_fu_2099_p2 = (add_ln703_345_fu_1970_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_305_fu_2104_p2 = (sub_ln703_286_fu_1989_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_306_fu_2109_p2 = (add_ln703_346_fu_1993_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_307_fu_2133_p2 = (sub_ln703_291_fu_2008_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_308_fu_2143_p2 = (add_ln703_348_fu_2017_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_309_fu_2148_p2 = (add_ln703_351_fu_2030_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_310_fu_2168_p2 = (sub_ln703_296_fu_2046_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_311_fu_2173_p2 = (add_ln703_352_fu_2051_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_312_fu_2409_p2 = (add_ln703_353_reg_5743 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_313_fu_2413_p2 = (sub_ln703_300_reg_5748 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_314_fu_2417_p2 = (add_ln703_354_reg_5753 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_315_fu_2188_p2 = (sub_ln703_301_fu_2085_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_316_fu_2421_p2 = (sub_ln703_302_reg_5758 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_317_fu_2425_p2 = (sub_ln703_304_reg_5763 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_318_fu_2203_p2 = (sub_ln703_306_fu_2109_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_319_fu_2208_p2 = (add_ln703_355_fu_2114_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_320_fu_2433_p2 = (add_ln703_359_reg_5768 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_321_fu_2218_p2 = (add_ln703_360_fu_2138_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_322_fu_2223_p2 = (sub_ln703_308_fu_2143_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_323_fu_2233_p2 = (add_ln703_362_fu_2158_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_324_fu_2238_p2 = (add_ln703_363_fu_2163_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_325_fu_2243_p2 = (sub_ln703_310_fu_2168_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_326_fu_2441_p2 = (sub_ln703_311_reg_5778 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_327_fu_2248_p2 = (add_ln703_364_fu_2178_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_328_fu_2253_p2 = (add_ln703_365_fu_2183_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_329_fu_2450_p2 = (sub_ln703_314_fu_2417_p2 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_330_fu_2455_p2 = (sub_ln703_316_fu_2421_p2 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_331_fu_2258_p2 = (add_ln703_366_fu_2193_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_332_fu_2273_p2 = (add_ln703_367_fu_2198_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_333_fu_2460_p2 = (sub_ln703_318_reg_5783 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_334_fu_2464_p2 = (add_ln703_368_fu_2429_p2 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_335_fu_2302_p2 = (add_ln703_369_fu_2213_p2 - data_20_V_read21_reg_4539_pp0_iter5_reg);

assign sub_ln703_336_fu_2469_p2 = (sub_ln703_321_reg_5788 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_337_fu_2473_p2 = (add_ln703_370_fu_2437_p2 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_338_fu_2478_p2 = (add_ln703_372_reg_5793 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_339_fu_2482_p2 = (sub_ln703_324_reg_5803 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_340_fu_2495_p2 = (sub_ln703_327_reg_5813 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_341_fu_2504_p2 = (add_ln703_373_fu_2445_p2 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_342_fu_2509_p2 = (sub_ln703_329_fu_2450_p2 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_343_fu_2312_p2 = (add_ln703_375_fu_2268_p2 - data_20_V_read21_reg_4539_pp0_iter5_reg);

assign sub_ln703_344_fu_2523_p2 = (add_ln703_377_reg_5833 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_345_fu_2532_p2 = (add_ln703_379_reg_5838 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_346_fu_2332_p2 = (add_ln703_380_fu_2297_p2 - data_20_V_read21_reg_4539_pp0_iter5_reg);

assign sub_ln703_347_fu_2536_p2 = (sub_ln703_335_reg_5843 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_348_fu_2545_p2 = (add_ln703_381_reg_5848 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_349_fu_2549_p2 = (sub_ln703_337_fu_2473_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_350_fu_2554_p2 = (sub_ln703_338_fu_2478_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_351_fu_2574_p2 = (sub_ln703_339_fu_2482_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_352_fu_2579_p2 = (add_ln703_382_fu_2486_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_353_fu_2584_p2 = (add_ln703_383_fu_2490_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_354_fu_2589_p2 = (sub_ln703_340_fu_2495_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_355_fu_2594_p2 = (add_ln703_385_fu_2499_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_356_fu_2603_p2 = (sub_ln703_341_fu_2504_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_357_fu_2608_p2 = (sub_ln703_342_fu_2509_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_358_fu_2613_p2 = (add_ln703_386_fu_2514_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_359_fu_2618_p2 = (add_ln703_387_fu_2518_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_360_fu_2627_p2 = (add_ln703_390_reg_5858 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_361_fu_2636_p2 = (add_ln703_391_fu_2527_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_362_fu_2641_p2 = (sub_ln703_346_reg_5863 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_363_fu_2660_p2 = (add_ln703_392_fu_2540_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_364_fu_2665_p2 = (sub_ln703_348_fu_2545_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_365_fu_2670_p2 = (sub_ln703_350_fu_2554_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_366_fu_2684_p2 = (add_ln703_396_fu_2568_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_367_fu_2689_p2 = (sub_ln703_351_fu_2574_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_368_fu_2694_p2 = (sub_ln703_352_fu_2579_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_369_fu_2699_p2 = (sub_ln703_353_fu_2584_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_370_fu_2714_p2 = (add_ln703_397_fu_2599_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_371_fu_2719_p2 = (add_ln703_400_reg_5868 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_372_fu_2985_p2 = (sub_ln703_356_reg_5921 - data_22_V_read23_reg_4483_pp0_iter7_reg);

assign sub_ln703_373_fu_2723_p2 = (sub_ln703_358_fu_2613_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_374_fu_2728_p2 = (sub_ln703_359_fu_2618_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_375_fu_2747_p2 = (add_ln703_401_fu_2623_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_376_fu_2752_p2 = (sub_ln703_360_fu_2627_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_377_fu_2989_p2 = (add_ln703_402_reg_5931 - data_22_V_read23_reg_4483_pp0_iter7_reg);

assign sub_ln703_378_fu_2776_p2 = (sub_ln703_362_fu_2641_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_379_fu_2781_p2 = (add_ln703_405_fu_2650_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_380_fu_2786_p2 = (add_ln703_406_fu_2655_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_381_fu_2791_p2 = (sub_ln703_363_fu_2660_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_382_fu_2796_p2 = (sub_ln703_364_fu_2665_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_383_fu_2801_p2 = (add_ln703_408_fu_2679_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_384_fu_2997_p2 = (sub_ln703_366_reg_5941 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_385_fu_2811_p2 = (sub_ln703_368_fu_2694_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_386_fu_2816_p2 = (add_ln703_409_fu_2704_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_387_fu_3005_p2 = (add_ln703_410_reg_5951 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_388_fu_2821_p2 = (add_ln703_413_reg_5873 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_389_fu_2839_p2 = (sub_ln703_371_fu_2719_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_390_fu_3009_p2 = (sub_ln703_372_fu_2985_p2 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_391_fu_2844_p2 = (add_ln703_415_reg_5878 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_392_fu_2848_p2 = (sub_ln703_373_fu_2723_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_393_fu_3018_p2 = (add_ln703_418_reg_5961 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_394_fu_3022_p2 = (sub_ln703_375_reg_5966 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_395_fu_2853_p2 = (sub_ln703_376_fu_2752_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_396_fu_2858_p2 = (add_ln703_420_fu_2761_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_397_fu_2863_p2 = (add_ln703_422_fu_2771_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_398_fu_3026_p2 = (sub_ln703_377_fu_2989_p2 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_399_fu_3031_p2 = (add_ln703_423_fu_2993_p2 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_400_fu_2868_p2 = (sub_ln703_378_fu_2776_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_401_fu_3040_p2 = (sub_ln703_381_reg_5976 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_402_fu_2878_p2 = (sub_ln703_382_fu_2796_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_403_fu_3044_p2 = (sub_ln703_384_fu_2997_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_404_fu_3049_p2 = (add_ln703_424_reg_5981 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_405_fu_3057_p2 = (add_ln703_425_fu_3001_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_406_fu_3062_p2 = (sub_ln703_386_reg_5991 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_407_fu_3066_p2 = (sub_ln703_387_fu_3005_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_408_fu_2893_p2 = (sub_ln703_388_fu_2821_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_409_fu_2898_p2 = (add_ln703_431_fu_2834_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_410_fu_3071_p2 = (sub_ln703_389_reg_5996 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_411_fu_2903_p2 = (sub_ln703_391_fu_2844_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_412_fu_3080_p2 = (sub_ln703_392_reg_6001 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_413_fu_3084_p2 = (add_ln703_432_fu_3014_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_414_fu_3089_p2 = (sub_ln703_393_fu_3018_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_415_fu_3094_p2 = (sub_ln703_394_fu_3022_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_416_fu_2923_p2 = (sub_ln703_396_fu_2858_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_417_fu_3103_p2 = (sub_ln703_399_fu_3031_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_418_fu_3108_p2 = (add_ln703_433_fu_3036_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_419_fu_3113_p2 = (add_ln703_434_reg_6011 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_420_fu_3117_p2 = (sub_ln703_401_fu_3040_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_421_fu_3126_p2 = (add_ln703_436_reg_6021 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_422_fu_3130_p2 = (sub_ln703_403_fu_3044_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_423_fu_3135_p2 = (sub_ln703_404_fu_3049_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_424_fu_3140_p2 = (add_ln703_437_fu_3053_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_425_fu_3145_p2 = (sub_ln703_406_fu_3062_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_426_fu_2938_p2 = (add_ln703_438_fu_2888_p2 - data_25_V_read26_reg_4391_pp0_iter6_reg);

assign sub_ln703_427_fu_3154_p2 = (sub_ln703_409_reg_6031 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_428_fu_3163_p2 = (add_ln703_439_fu_3075_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_429_fu_3177_p2 = (sub_ln703_411_reg_6036 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_430_fu_3181_p2 = (add_ln703_442_reg_6041 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_431_fu_3185_p2 = (sub_ln703_412_fu_3080_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_432_fu_3190_p2 = (sub_ln703_416_reg_6046 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_433_fu_3194_p2 = (add_ln703_443_fu_3099_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_434_fu_3199_p2 = (sub_ln703_417_fu_3103_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_435_fu_3204_p2 = (add_ln703_444_reg_6051 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_436_fu_3208_p2 = (sub_ln703_418_fu_3108_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_437_fu_3213_p2 = (sub_ln703_419_fu_3113_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_438_fu_3223_p2 = (add_ln703_445_fu_3122_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_439_fu_3228_p2 = (add_ln703_447_reg_6056 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_440_fu_3247_p2 = (sub_ln703_425_fu_3145_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_441_fu_3252_p2 = (sub_ln703_426_reg_6061 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_442_fu_3256_p2 = (add_ln703_448_fu_3150_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_443_fu_3261_p2 = (sub_ln703_427_fu_3154_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_444_fu_3266_p2 = (add_ln703_449_fu_3158_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_445_fu_3271_p2 = (add_ln703_452_fu_3172_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_446_fu_3276_p2 = (sub_ln703_429_fu_3177_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_447_fu_3298_p2 = (sub_ln703_432_fu_3190_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_448_fu_3308_p2 = (sub_ln703_436_fu_3208_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_449_fu_3313_p2 = (sub_ln703_437_fu_3213_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_450_fu_3318_p2 = (add_ln703_453_fu_3218_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_451_fu_3343_p2 = (add_ln703_454_fu_3232_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_452_fu_3348_p2 = (add_ln703_456_fu_3241_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_453_fu_3353_p2 = (sub_ln703_440_fu_3247_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_454_fu_3368_p2 = (sub_ln703_441_fu_3252_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_455_fu_3373_p2 = (sub_ln703_444_fu_3266_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_456_fu_3388_p2 = (add_ln703_457_fu_3281_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_457_fu_3393_p2 = (add_ln703_458_fu_3286_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_458_fu_3408_p2 = (add_ln703_459_fu_3292_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_459_fu_3418_p2 = (add_ln703_460_fu_3303_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_460_fu_3535_p2 = (sub_ln703_450_reg_6123 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_461_fu_3438_p2 = (add_ln703_461_fu_3323_p2 - data_28_V_read_7_reg_4313_pp0_iter7_reg);

assign sub_ln703_462_fu_3539_p2 = (add_ln703_463_reg_6128 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_463_fu_3543_p2 = (add_ln703_464_reg_6133 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_464_fu_3547_p2 = (add_ln703_465_reg_6138 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_465_fu_3551_p2 = (sub_ln703_451_reg_6143 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_466_fu_3563_p2 = (add_ln703_467_reg_6158 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_467_fu_3567_p2 = (sub_ln703_454_reg_6163 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_468_fu_3575_p2 = (add_ln703_468_reg_6173 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_469_fu_3463_p2 = (add_ln703_469_fu_3383_p2 - data_28_V_read_7_reg_4313_pp0_iter7_reg);

assign sub_ln703_470_fu_3579_p2 = (sub_ln703_456_reg_6178 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_471_fu_3583_p2 = (sub_ln703_457_reg_6183 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_472_fu_3587_p2 = (add_ln703_471_reg_6188 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_473_fu_3591_p2 = (sub_ln703_458_reg_6193 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_474_fu_3482_p2 = (add_ln703_472_fu_3413_p2 - data_28_V_read_7_reg_4313_pp0_iter7_reg);

assign sub_ln703_475_fu_3599_p2 = (sub_ln703_459_reg_6198 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_476_fu_3603_p2 = (add_ln703_475_reg_6203 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_477_fu_3607_p2 = (add_ln703_476_fu_3531_p2 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_478_fu_3612_p2 = (add_ln703_480_reg_6072_pp0_iter8_reg - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_479_fu_3621_p2 = (sub_ln703_462_fu_3539_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_480_fu_3626_p2 = (sub_ln703_463_fu_3543_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_481_fu_3636_p2 = (add_ln703_483_reg_6213 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_482_fu_3640_p2 = (sub_ln703_465_fu_3551_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_483_fu_3645_p2 = (add_ln703_484_fu_3555_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_484_fu_3650_p2 = (add_ln703_485_fu_3559_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_485_fu_3660_p2 = (sub_ln703_467_fu_3567_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_486_fu_3507_p2 = (add_ln703_486_fu_3453_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_487_fu_3512_p2 = (add_ln703_487_fu_3458_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_488_fu_3665_p2 = (add_ln703_488_fu_3571_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_489_fu_3670_p2 = (sub_ln703_468_fu_3575_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_490_fu_3675_p2 = (sub_ln703_469_reg_6218 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_491_fu_3517_p2 = (add_ln703_490_fu_3473_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_492_fu_3679_p2 = (sub_ln703_470_fu_3579_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_493_fu_3684_p2 = (sub_ln703_471_fu_3583_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_494_fu_3689_p2 = (sub_ln703_472_fu_3587_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_495_fu_3694_p2 = (sub_ln703_473_fu_3591_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_496_fu_3699_p2 = (add_ln703_493_fu_3595_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_497_fu_3704_p2 = (sub_ln703_474_reg_6229 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_498_fu_3718_p2 = (sub_ln703_477_fu_3607_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_499_fu_3723_p2 = (sub_ln703_478_fu_3612_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_500_fu_3522_p2 = (add_ln703_495_fu_3492_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_501_fu_3728_p2 = (add_ln703_497_reg_6239 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_502_fu_3732_p2 = (add_ln703_498_fu_3616_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_503_fu_3737_p2 = (sub_ln703_479_fu_3621_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_504_fu_3742_p2 = (sub_ln703_480_fu_3626_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_505_fu_3747_p2 = (add_ln703_499_fu_3631_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_506_fu_3752_p2 = (sub_ln703_482_fu_3640_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_507_fu_3762_p2 = (sub_ln703_484_fu_3650_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_508_fu_3767_p2 = (add_ln703_500_fu_3655_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_509_fu_3772_p2 = (sub_ln703_485_fu_3660_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_510_fu_3781_p2 = (sub_ln703_487_reg_6249 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_511_fu_3790_p2 = (sub_ln703_489_fu_3670_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_512_fu_3804_p2 = (sub_ln703_493_fu_3684_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_513_fu_3809_p2 = (sub_ln703_494_fu_3689_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_514_fu_3814_p2 = (sub_ln703_495_fu_3694_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_515_fu_3819_p2 = (sub_ln703_496_fu_3699_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_516_fu_3824_p2 = (add_ln703_501_fu_3708_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_517_fu_3829_p2 = (add_ln703_502_fu_3713_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_518_fu_3834_p2 = (sub_ln703_499_fu_3723_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_519_fu_3839_p2 = (sub_ln703_500_reg_6259 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_73_fu_286_p2 = (data_0_V_read_int_reg - data_1_V_read_int_reg);

assign sub_ln703_74_fu_292_p2 = (sub_ln703_reg_5046 - data_2_V_read_9_reg_5035);

assign sub_ln703_75_fu_296_p2 = (add_ln703_reg_5052 - data_2_V_read_9_reg_5035);

assign sub_ln703_76_fu_300_p2 = (sub_ln703_73_reg_5059 - data_2_V_read_9_reg_5035);

assign sub_ln703_77_fu_308_p2 = (data_2_V_read_9_reg_5035 - add_ln703_reg_5052);

assign sub_ln703_78_fu_361_p2 = (sub_ln703_76_reg_5071_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_79_fu_337_p2 = (sub_ln703_77_reg_5084 - data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign sub_ln703_80_fu_365_p2 = (add_ln703_201_reg_5090_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_81_fu_369_p2 = (add_ln703_202_reg_5096_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_82_fu_373_p2 = (data_3_V_read_9_reg_5019_pp0_iter2_reg - add_ln703_200_reg_5077_pp0_iter2_reg);

assign sub_ln703_83_fu_377_p2 = (add_ln703_200_reg_5077_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_84_fu_381_p2 = (sub_ln703_74_reg_5065_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_85_fu_385_p2 = (add_ln703_203_reg_5113 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_86_fu_389_p2 = (add_ln703_204_reg_5101_pp0_iter2_reg - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_87_fu_393_p2 = (sub_ln703_78_fu_361_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_88_fu_398_p2 = (data_4_V_read_9_reg_4998_pp0_iter2_reg - add_ln703_205_reg_5119);

assign sub_ln703_89_fu_402_p2 = (sub_ln703_79_reg_5125 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_90_fu_406_p2 = (sub_ln703_80_fu_365_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_91_fu_411_p2 = (sub_ln703_81_fu_369_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_92_fu_437_p2 = (sub_ln703_84_fu_381_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_93_fu_442_p2 = (add_ln703_206_reg_5131 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_94_fu_446_p2 = (sub_ln703_86_fu_389_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_95_fu_451_p2 = (sub_ln703_87_fu_393_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_96_fu_456_p2 = (sub_ln703_88_fu_398_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_97_fu_609_p2 = (sub_ln703_91_reg_5172 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_98_fu_466_p2 = (add_ln703_208_reg_5137 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_99_fu_613_p2 = (data_5_V_read_8_reg_4969_pp0_iter3_reg - add_ln703_209_reg_5178);

assign sub_ln703_fu_274_p2 = (data_1_V_read_int_reg - data_0_V_read_int_reg);

endmodule //dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        data_32_V_read,
        data_33_V_read,
        data_34_V_read,
        data_35_V_read,
        data_36_V_read,
        data_37_V_read,
        data_38_V_read,
        data_39_V_read,
        data_40_V_read,
        data_41_V_read,
        data_42_V_read,
        data_43_V_read,
        data_44_V_read,
        data_45_V_read,
        data_46_V_read,
        data_47_V_read,
        data_48_V_read,
        data_49_V_read,
        data_50_V_read,
        data_51_V_read,
        data_52_V_read,
        data_53_V_read,
        data_54_V_read,
        data_55_V_read,
        data_56_V_read,
        data_57_V_read,
        data_58_V_read,
        data_59_V_read,
        data_60_V_read,
        data_61_V_read,
        data_62_V_read,
        data_63_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
input  [15:0] data_32_V_read;
input  [15:0] data_33_V_read;
input  [15:0] data_34_V_read;
input  [15:0] data_35_V_read;
input  [15:0] data_36_V_read;
input  [15:0] data_37_V_read;
input  [15:0] data_38_V_read;
input  [15:0] data_39_V_read;
input  [15:0] data_40_V_read;
input  [15:0] data_41_V_read;
input  [15:0] data_42_V_read;
input  [15:0] data_43_V_read;
input  [15:0] data_44_V_read;
input  [15:0] data_45_V_read;
input  [15:0] data_46_V_read;
input  [15:0] data_47_V_read;
input  [15:0] data_48_V_read;
input  [15:0] data_49_V_read;
input  [15:0] data_50_V_read;
input  [15:0] data_51_V_read;
input  [15:0] data_52_V_read;
input  [15:0] data_53_V_read;
input  [15:0] data_54_V_read;
input  [15:0] data_55_V_read;
input  [15:0] data_56_V_read;
input  [15:0] data_57_V_read;
input  [15:0] data_58_V_read;
input  [15:0] data_59_V_read;
input  [15:0] data_60_V_read;
input  [15:0] data_61_V_read;
input  [15:0] data_62_V_read;
input  [15:0] data_63_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;

reg   [15:0] data_63_V_read_3_reg_8620;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter1_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter2_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter3_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter4_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter5_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter6_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter7_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter8_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter9_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter10_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter11_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter12_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter13_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter14_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter15_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter16_reg;
reg   [15:0] data_62_V_read_3_reg_8645;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter1_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter2_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter3_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter4_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter5_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter6_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter7_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter8_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter9_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter10_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter11_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter12_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter13_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter14_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter15_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter16_reg;
reg   [15:0] data_61_V_read62_reg_8663;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter1_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter2_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter3_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter4_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter5_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter6_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter7_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter8_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter9_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter10_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter11_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter12_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter13_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter14_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter15_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter16_reg;
reg   [15:0] data_60_V_read61_reg_8691;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter1_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter2_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter3_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter4_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter5_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter6_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter7_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter8_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter9_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter10_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter11_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter12_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter13_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter14_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter15_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter16_reg;
reg   [15:0] data_59_V_read_3_reg_8724;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter1_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter2_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter3_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter4_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter5_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter6_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter7_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter8_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter9_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter10_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter11_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter12_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter13_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter14_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter15_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter16_reg;
reg   [15:0] data_58_V_read_3_reg_8756;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter1_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter2_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter3_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter4_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter5_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter6_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter7_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter8_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter9_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter10_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter11_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter12_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter13_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter14_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter15_reg;
reg   [15:0] data_57_V_read_3_reg_8786;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter1_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter2_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter3_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter4_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter5_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter6_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter7_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter8_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter9_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter10_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter11_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter12_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter13_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter14_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter15_reg;
reg   [15:0] data_56_V_read_3_reg_8814;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter1_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter2_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter3_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter4_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter5_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter6_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter7_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter8_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter9_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter10_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter11_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter12_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter13_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter14_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter15_reg;
reg   [15:0] data_55_V_read_3_reg_8844;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter1_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter2_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter3_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter4_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter5_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter6_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter7_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter8_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter9_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter10_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter11_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter12_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter13_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter14_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter15_reg;
reg   [15:0] data_54_V_read_3_reg_8873;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter1_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter2_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter3_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter4_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter5_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter6_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter7_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter8_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter9_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter10_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter11_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter12_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter13_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter14_reg;
reg   [15:0] data_53_V_read_3_reg_8899;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter1_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter2_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter3_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter4_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter5_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter6_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter7_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter8_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter9_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter10_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter11_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter12_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter13_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter14_reg;
reg   [15:0] data_52_V_read_3_reg_8928;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter1_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter2_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter3_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter4_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter5_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter6_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter7_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter8_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter9_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter10_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter11_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter12_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter13_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter14_reg;
reg   [15:0] data_51_V_read52_reg_8956;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter1_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter2_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter3_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter4_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter5_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter6_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter7_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter8_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter9_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter10_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter11_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter12_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter13_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter14_reg;
reg   [15:0] data_50_V_read51_reg_8984;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter1_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter2_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter3_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter4_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter5_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter6_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter7_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter8_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter9_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter10_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter11_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter12_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter13_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter14_reg;
reg   [15:0] data_49_V_read_3_reg_9012;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter1_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter2_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter3_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter4_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter5_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter6_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter7_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter8_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter9_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter10_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter11_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter12_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter13_reg;
reg   [15:0] data_48_V_read_3_reg_9040;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter1_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter2_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter3_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter4_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter5_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter6_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter7_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter8_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter9_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter10_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter11_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter12_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter13_reg;
reg   [15:0] data_47_V_read_3_reg_9066;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter1_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter2_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter3_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter4_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter5_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter6_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter7_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter8_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter9_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter10_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter11_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter12_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter13_reg;
reg   [15:0] data_46_V_read_3_reg_9094;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter1_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter2_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter3_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter4_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter5_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter6_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter7_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter8_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter9_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter10_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter11_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter12_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter13_reg;
reg   [15:0] data_45_V_read_3_reg_9125;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter1_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter2_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter3_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter4_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter5_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter6_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter7_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter8_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter9_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter10_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter11_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter12_reg;
reg   [15:0] data_44_V_read_3_reg_9154;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter1_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter2_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter3_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter4_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter5_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter6_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter7_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter8_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter9_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter10_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter11_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter12_reg;
reg   [15:0] data_43_V_read_3_reg_9184;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter1_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter2_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter3_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter4_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter5_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter6_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter7_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter8_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter9_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter10_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter11_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter12_reg;
reg   [15:0] data_42_V_read_3_reg_9212;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter1_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter2_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter3_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter4_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter5_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter6_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter7_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter8_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter9_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter10_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter11_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter12_reg;
reg   [15:0] data_41_V_read42_reg_9242;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter1_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter2_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter3_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter4_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter5_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter6_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter7_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter8_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter9_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter10_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter11_reg;
reg   [15:0] data_40_V_read41_reg_9272;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter1_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter2_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter3_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter4_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter5_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter6_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter7_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter8_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter9_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter10_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter11_reg;
reg   [15:0] data_39_V_read_3_reg_9301;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter1_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter2_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter3_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter4_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter5_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter6_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter7_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter8_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter9_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter10_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter11_reg;
reg   [15:0] data_38_V_read_3_reg_9328;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter1_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter2_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter3_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter4_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter5_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter6_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter7_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter8_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter9_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter10_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter11_reg;
reg   [15:0] data_37_V_read_3_reg_9353;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter1_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter2_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter3_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter4_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter5_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter6_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter7_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter8_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter9_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter10_reg;
reg   [15:0] data_36_V_read_3_reg_9383;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter1_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter2_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter3_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter4_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter5_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter6_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter7_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter8_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter9_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter10_reg;
reg   [15:0] data_35_V_read_3_reg_9410;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter1_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter2_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter3_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter4_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter5_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter6_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter7_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter8_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter9_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter10_reg;
reg   [15:0] data_34_V_read_3_reg_9434;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter1_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter2_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter3_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter4_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter5_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter6_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter7_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter8_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter9_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter10_reg;
reg   [15:0] data_33_V_read_3_reg_9463;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter1_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter2_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter3_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter4_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter5_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter6_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter7_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter8_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter9_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter10_reg;
reg   [15:0] data_32_V_read_3_reg_9492;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter1_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter2_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter3_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter4_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter5_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter6_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter7_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter8_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter9_reg;
reg   [15:0] data_31_V_read32_reg_9521;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter1_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter2_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter3_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter4_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter5_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter6_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter7_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter8_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter9_reg;
reg   [15:0] data_30_V_read31_reg_9549;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter1_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter2_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter3_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter4_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter5_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter6_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter7_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter8_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter9_reg;
reg   [15:0] data_29_V_read_8_reg_9573;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter1_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter2_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter3_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter4_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter5_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter6_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter7_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter8_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter9_reg;
reg   [15:0] data_28_V_read_8_reg_9598;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter1_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter2_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter3_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter4_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter5_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter6_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter7_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter8_reg;
reg   [15:0] data_27_V_read28_reg_9625;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter1_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter2_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter3_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter4_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter5_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter6_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter7_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter8_reg;
reg   [15:0] data_26_V_read27_reg_9652;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter1_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter2_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter3_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter4_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter5_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter6_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter7_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter8_reg;
reg   [15:0] data_25_V_read26_reg_9677;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter1_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter2_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter3_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter4_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter5_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter6_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter7_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter8_reg;
reg   [15:0] data_24_V_read25_reg_9704;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter1_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter2_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter3_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter4_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter5_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter6_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter7_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter8_reg;
reg   [15:0] data_23_V_read24_reg_9730;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter1_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter2_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter3_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter4_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter5_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter6_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter7_reg;
reg   [15:0] data_22_V_read23_reg_9756;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter1_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter2_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter3_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter5_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter6_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter7_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter8_reg;
reg   [15:0] data_21_V_read22_reg_9784;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter1_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter2_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter3_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter4_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter5_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter6_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter7_reg;
reg   [15:0] data_20_V_read21_reg_9814;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter1_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter2_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter3_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter4_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter5_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter6_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter7_reg;
reg   [15:0] data_19_V_read_8_reg_9845;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter1_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter2_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter3_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter4_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter5_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter6_reg;
reg   [15:0] data_18_V_read_8_reg_9874;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter1_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter2_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter3_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter4_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter5_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter6_reg;
reg   [15:0] data_17_V_read18_reg_9904;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter1_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter2_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter3_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter4_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter5_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter6_reg;
reg   [15:0] data_16_V_read17_reg_9935;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter1_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter2_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter3_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter4_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter5_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter6_reg;
reg   [15:0] data_15_V_read16_reg_9962;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter1_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter2_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter3_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter4_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter5_reg;
reg   [15:0] data_14_V_read15_reg_9987;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter1_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter2_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter3_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter4_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter5_reg;
reg   [15:0] data_13_V_read14_reg_10015;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter1_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter2_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter3_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter4_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter5_reg;
reg   [15:0] data_12_V_read13_reg_10045;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter1_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter2_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter3_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter4_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter5_reg;
reg   [15:0] data_11_V_read12_reg_10075;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter1_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter2_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter3_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter4_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter5_reg;
reg   [15:0] data_10_V_read11_reg_10105;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter1_reg;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter2_reg;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter3_reg;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter4_reg;
reg   [15:0] data_9_V_read_8_reg_10136;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter1_reg;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter2_reg;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter3_reg;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter4_reg;
reg   [15:0] data_8_V_read_8_reg_10164;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter1_reg;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter2_reg;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter3_reg;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter4_reg;
reg   [15:0] data_7_V_read_9_reg_10191;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter1_reg;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter2_reg;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter3_reg;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter4_reg;
reg   [15:0] data_6_V_read_9_reg_10218;
reg   [15:0] data_6_V_read_9_reg_10218_pp0_iter1_reg;
reg   [15:0] data_6_V_read_9_reg_10218_pp0_iter2_reg;
reg   [15:0] data_6_V_read_9_reg_10218_pp0_iter3_reg;
reg   [15:0] data_5_V_read_9_reg_10245;
reg   [15:0] data_5_V_read_9_reg_10245_pp0_iter1_reg;
reg   [15:0] data_5_V_read_9_reg_10245_pp0_iter2_reg;
reg   [15:0] data_5_V_read_9_reg_10245_pp0_iter3_reg;
reg   [15:0] data_4_V_read_10_reg_10273;
reg   [15:0] data_4_V_read_10_reg_10273_pp0_iter1_reg;
reg   [15:0] data_4_V_read_10_reg_10273_pp0_iter2_reg;
reg   [15:0] data_4_V_read_10_reg_10273_pp0_iter3_reg;
reg   [15:0] data_3_V_read_10_reg_10295;
reg   [15:0] data_3_V_read_10_reg_10295_pp0_iter1_reg;
reg   [15:0] data_3_V_read_10_reg_10295_pp0_iter2_reg;
reg   [15:0] data_2_V_read_10_reg_10312;
reg   [15:0] data_2_V_read_10_reg_10312_pp0_iter1_reg;
reg   [15:0] data_1_V_read_10_reg_10323;
reg   [15:0] data_0_V_read_10_reg_10329;
wire   [15:0] add_ln703_fu_530_p2;
reg   [15:0] add_ln703_reg_10335;
reg   [15:0] add_ln703_reg_10335_pp0_iter1_reg;
wire   [15:0] sub_ln703_fu_536_p2;
reg   [15:0] sub_ln703_reg_10342;
wire   [15:0] sub_ln703_1_fu_540_p2;
reg   [15:0] sub_ln703_1_reg_10348;
wire   [15:0] add_ln703_131_fu_544_p2;
reg   [15:0] add_ln703_131_reg_10354;
reg   [15:0] add_ln703_131_reg_10354_pp0_iter2_reg;
wire   [15:0] sub_ln703_4_fu_548_p2;
reg   [15:0] sub_ln703_4_reg_10361;
reg   [15:0] sub_ln703_4_reg_10361_pp0_iter2_reg;
wire   [15:0] sub_ln703_2_fu_552_p2;
reg   [15:0] sub_ln703_2_reg_10367;
wire   [15:0] add_ln703_130_fu_556_p2;
reg   [15:0] add_ln703_130_reg_10373;
wire   [15:0] sub_ln703_3_fu_560_p2;
reg   [15:0] sub_ln703_3_reg_10379;
wire   [15:0] add_ln703_134_fu_568_p2;
reg   [15:0] add_ln703_134_reg_10385;
wire   [15:0] sub_ln703_8_fu_572_p2;
reg   [15:0] sub_ln703_8_reg_10392;
wire   [15:0] sub_ln703_11_fu_576_p2;
reg   [15:0] sub_ln703_11_reg_10398;
reg   [15:0] sub_ln703_11_reg_10398_pp0_iter3_reg;
wire   [15:0] add_ln703_144_fu_589_p2;
reg   [15:0] add_ln703_144_reg_10403;
reg   [15:0] add_ln703_144_reg_10403_pp0_iter3_reg;
wire   [15:0] sub_ln703_6_fu_595_p2;
reg   [15:0] sub_ln703_6_reg_10408;
wire   [15:0] add_ln703_132_fu_599_p2;
reg   [15:0] add_ln703_132_reg_10414;
wire   [15:0] sub_ln703_10_fu_615_p2;
reg   [15:0] sub_ln703_10_reg_10420;
wire   [15:0] add_ln703_135_fu_619_p2;
reg   [15:0] add_ln703_135_reg_10425;
wire   [15:0] sub_ln703_15_fu_631_p2;
reg   [15:0] sub_ln703_15_reg_10430;
wire   [15:0] sub_ln703_16_fu_640_p2;
reg   [15:0] sub_ln703_16_reg_10436;
wire   [15:0] add_ln703_140_fu_644_p2;
reg   [15:0] add_ln703_140_reg_10442;
wire   [15:0] add_ln703_141_fu_649_p2;
reg   [15:0] add_ln703_141_reg_10447;
wire   [15:0] sub_ln703_17_fu_653_p2;
reg   [15:0] sub_ln703_17_reg_10453;
wire   [15:0] sub_ln703_18_fu_658_p2;
reg   [15:0] sub_ln703_18_reg_10459;
wire   [15:0] sub_ln703_20_fu_662_p2;
reg   [15:0] sub_ln703_20_reg_10465;
wire   [15:0] sub_ln703_23_fu_666_p2;
reg   [15:0] sub_ln703_23_reg_10471;
wire   [15:0] sub_ln703_28_fu_671_p2;
reg   [15:0] sub_ln703_28_reg_10476;
wire   [15:0] add_ln703_158_fu_676_p2;
reg   [15:0] add_ln703_158_reg_10482;
wire   [15:0] add_ln703_161_fu_681_p2;
reg   [15:0] add_ln703_161_reg_10487;
wire   [15:0] add_ln703_179_fu_685_p2;
reg   [15:0] add_ln703_179_reg_10495;
wire   [15:0] add_ln703_153_fu_809_p2;
reg   [15:0] add_ln703_153_reg_10503;
wire   [15:0] sub_ln703_38_fu_814_p2;
reg   [15:0] sub_ln703_38_reg_10508;
wire   [15:0] sub_ln703_39_fu_819_p2;
reg   [15:0] sub_ln703_39_reg_10513;
wire   [15:0] sub_ln703_40_fu_824_p2;
reg   [15:0] sub_ln703_40_reg_10519;
wire   [15:0] sub_ln703_43_fu_838_p2;
reg   [15:0] sub_ln703_43_reg_10524;
wire   [15:0] add_ln703_157_fu_892_p2;
reg   [15:0] add_ln703_157_reg_10529;
wire   [15:0] sub_ln703_53_fu_912_p2;
reg   [15:0] sub_ln703_53_reg_10534;
wire   [15:0] add_ln703_162_fu_917_p2;
reg   [15:0] add_ln703_162_reg_10539;
wire   [15:0] sub_ln703_58_fu_922_p2;
reg   [15:0] sub_ln703_58_reg_10545;
wire   [15:0] sub_ln703_62_fu_942_p2;
reg   [15:0] sub_ln703_62_reg_10550;
wire   [15:0] sub_ln703_63_fu_947_p2;
reg   [15:0] sub_ln703_63_reg_10555;
wire   [15:0] sub_ln703_64_fu_957_p2;
reg   [15:0] sub_ln703_64_reg_10560;
wire   [15:0] add_ln703_170_fu_972_p2;
reg   [15:0] add_ln703_170_reg_10566;
wire   [15:0] add_ln703_171_fu_977_p2;
reg   [15:0] add_ln703_171_reg_10571;
wire   [15:0] add_ln703_173_fu_982_p2;
reg   [15:0] add_ln703_173_reg_10576;
wire   [15:0] sub_ln703_66_fu_987_p2;
reg   [15:0] sub_ln703_66_reg_10581;
wire   [15:0] sub_ln703_70_fu_992_p2;
reg   [15:0] sub_ln703_70_reg_10586;
wire   [15:0] add_ln703_177_fu_997_p2;
reg   [15:0] add_ln703_177_reg_10591;
wire   [15:0] sub_ln703_71_fu_1002_p2;
reg   [15:0] sub_ln703_71_reg_10596;
wire   [15:0] add_ln703_181_fu_1015_p2;
reg   [15:0] add_ln703_181_reg_10601;
wire   [15:0] add_ln703_183_fu_1021_p2;
reg   [15:0] add_ln703_183_reg_10606;
wire   [15:0] sub_ln703_73_fu_1026_p2;
reg   [15:0] sub_ln703_73_reg_10611;
wire   [15:0] sub_ln703_75_fu_1031_p2;
reg   [15:0] sub_ln703_75_reg_10616;
wire   [15:0] add_ln703_186_fu_1036_p2;
reg   [15:0] add_ln703_186_reg_10621;
wire   [15:0] add_ln703_192_fu_1050_p2;
reg   [15:0] add_ln703_192_reg_10626;
wire   [15:0] sub_ln703_92_fu_1054_p2;
reg   [15:0] sub_ln703_92_reg_10636;
wire   [15:0] add_ln703_204_fu_1059_p2;
reg   [15:0] add_ln703_204_reg_10641;
wire   [15:0] add_ln703_209_fu_1064_p2;
reg   [15:0] add_ln703_209_reg_10646;
wire   [15:0] add_ln703_213_fu_1068_p2;
reg   [15:0] add_ln703_213_reg_10653;
wire   [15:0] add_ln703_223_fu_1073_p2;
reg   [15:0] add_ln703_223_reg_10658;
wire   [15:0] add_ln703_252_fu_1077_p2;
reg   [15:0] add_ln703_252_reg_10665;
reg   [15:0] add_ln703_252_reg_10665_pp0_iter5_reg;
wire   [15:0] add_ln703_254_fu_1081_p2;
reg   [15:0] add_ln703_254_reg_10672;
wire   [15:0] sub_ln703_96_fu_1294_p2;
reg   [15:0] sub_ln703_96_reg_10677;
wire   [15:0] add_ln703_207_fu_1299_p2;
reg   [15:0] add_ln703_207_reg_10682;
wire   [15:0] add_ln703_208_fu_1309_p2;
reg   [15:0] add_ln703_208_reg_10687;
wire   [15:0] add_ln703_210_fu_1314_p2;
reg   [15:0] add_ln703_210_reg_10692;
wire   [15:0] sub_ln703_98_fu_1319_p2;
reg   [15:0] sub_ln703_98_reg_10697;
wire   [15:0] add_ln703_216_fu_1358_p2;
reg   [15:0] add_ln703_216_reg_10702;
wire   [15:0] sub_ln703_106_fu_1378_p2;
reg   [15:0] sub_ln703_106_reg_10707;
wire   [15:0] sub_ln703_107_fu_1383_p2;
reg   [15:0] sub_ln703_107_reg_10712;
wire   [15:0] sub_ln703_108_fu_1388_p2;
reg   [15:0] sub_ln703_108_reg_10717;
wire   [15:0] sub_ln703_109_fu_1407_p2;
reg   [15:0] sub_ln703_109_reg_10722;
wire   [15:0] sub_ln703_115_fu_1432_p2;
reg   [15:0] sub_ln703_115_reg_10727;
wire   [15:0] add_ln703_224_fu_1437_p2;
reg   [15:0] add_ln703_224_reg_10732;
wire   [15:0] add_ln703_226_fu_1457_p2;
reg   [15:0] add_ln703_226_reg_10737;
wire   [15:0] sub_ln703_122_fu_1462_p2;
reg   [15:0] sub_ln703_122_reg_10742;
wire   [15:0] sub_ln703_123_fu_1467_p2;
reg   [15:0] sub_ln703_123_reg_10747;
wire   [15:0] add_ln703_227_fu_1472_p2;
reg   [15:0] add_ln703_227_reg_10752;
wire   [15:0] sub_ln703_125_fu_1482_p2;
reg   [15:0] sub_ln703_125_reg_10757;
wire   [15:0] sub_ln703_128_fu_1496_p2;
reg   [15:0] sub_ln703_128_reg_10762;
wire   [15:0] add_ln703_233_fu_1501_p2;
reg   [15:0] add_ln703_233_reg_10767;
wire   [15:0] add_ln703_236_fu_1511_p2;
reg   [15:0] add_ln703_236_reg_10772;
wire   [15:0] add_ln703_238_fu_1520_p2;
reg   [15:0] add_ln703_238_reg_10777;
wire   [15:0] sub_ln703_133_fu_1532_p2;
reg   [15:0] sub_ln703_133_reg_10782;
wire   [15:0] sub_ln703_137_fu_1548_p2;
reg   [15:0] sub_ln703_137_reg_10787;
wire   [15:0] sub_ln703_141_fu_1553_p2;
reg   [15:0] sub_ln703_141_reg_10792;
wire   [15:0] sub_ln703_142_fu_1558_p2;
reg   [15:0] sub_ln703_142_reg_10797;
wire   [15:0] add_ln703_247_fu_1563_p2;
reg   [15:0] add_ln703_247_reg_10802;
wire   [15:0] add_ln703_250_fu_1574_p2;
reg   [15:0] add_ln703_250_reg_10807;
wire   [15:0] sub_ln703_146_fu_1580_p2;
reg   [15:0] sub_ln703_146_reg_10812;
wire   [15:0] add_ln703_260_fu_1593_p2;
reg   [15:0] add_ln703_260_reg_10817;
wire   [15:0] sub_ln703_152_fu_1599_p2;
reg   [15:0] sub_ln703_152_reg_10822;
wire   [15:0] add_ln703_262_fu_1604_p2;
reg   [15:0] add_ln703_262_reg_10827;
wire   [15:0] sub_ln703_154_fu_1609_p2;
reg   [15:0] sub_ln703_154_reg_10832;
wire   [15:0] add_ln703_265_fu_1614_p2;
reg   [15:0] add_ln703_265_reg_10837;
wire   [15:0] add_ln703_280_fu_1618_p2;
reg   [15:0] add_ln703_280_reg_10846;
wire   [15:0] add_ln703_326_fu_1622_p2;
reg   [15:0] add_ln703_326_reg_10855;
reg   [15:0] add_ln703_326_reg_10855_pp0_iter6_reg;
wire   [15:0] sub_ln703_166_fu_1834_p2;
reg   [15:0] sub_ln703_166_reg_10863;
wire   [15:0] sub_ln703_183_fu_1959_p2;
reg   [15:0] sub_ln703_183_reg_10868;
wire   [15:0] add_ln703_283_fu_1979_p2;
reg   [15:0] add_ln703_283_reg_10873;
wire   [15:0] sub_ln703_184_fu_1984_p2;
reg   [15:0] sub_ln703_184_reg_10878;
wire   [15:0] sub_ln703_186_fu_1994_p2;
reg   [15:0] sub_ln703_186_reg_10883;
wire   [15:0] add_ln703_285_fu_2009_p2;
reg   [15:0] add_ln703_285_reg_10888;
wire   [15:0] sub_ln703_191_fu_2029_p2;
reg   [15:0] sub_ln703_191_reg_10893;
wire   [15:0] add_ln703_289_fu_2034_p2;
reg   [15:0] add_ln703_289_reg_10898;
wire   [15:0] add_ln703_290_fu_2039_p2;
reg   [15:0] add_ln703_290_reg_10903;
wire   [15:0] sub_ln703_194_fu_2054_p2;
reg   [15:0] sub_ln703_194_reg_10908;
wire   [15:0] sub_ln703_196_fu_2074_p2;
reg   [15:0] sub_ln703_196_reg_10913;
wire   [15:0] add_ln703_294_fu_2084_p2;
reg   [15:0] add_ln703_294_reg_10918;
wire   [15:0] add_ln703_295_fu_2089_p2;
reg   [15:0] add_ln703_295_reg_10923;
wire   [15:0] add_ln703_300_fu_2093_p2;
reg   [15:0] add_ln703_300_reg_10930;
wire   [15:0] sub_ln703_198_fu_2099_p2;
reg   [15:0] sub_ln703_198_reg_10935;
wire   [15:0] add_ln703_303_fu_2104_p2;
reg   [15:0] add_ln703_303_reg_10940;
wire   [15:0] add_ln703_304_fu_2110_p2;
reg   [15:0] add_ln703_304_reg_10945;
wire   [15:0] sub_ln703_200_fu_2115_p2;
reg   [15:0] sub_ln703_200_reg_10950;
wire   [15:0] sub_ln703_202_fu_2120_p2;
reg   [15:0] sub_ln703_202_reg_10955;
wire   [15:0] add_ln703_307_fu_2125_p2;
reg   [15:0] add_ln703_307_reg_10960;
wire   [15:0] sub_ln703_203_fu_2131_p2;
reg   [15:0] sub_ln703_203_reg_10965;
wire   [15:0] add_ln703_309_fu_2136_p2;
reg   [15:0] add_ln703_309_reg_10970;
wire   [15:0] sub_ln703_204_fu_2142_p2;
reg   [15:0] sub_ln703_204_reg_10975;
wire   [15:0] add_ln703_310_fu_2147_p2;
reg   [15:0] add_ln703_310_reg_10980;
wire   [15:0] sub_ln703_208_fu_2152_p2;
reg   [15:0] sub_ln703_208_reg_10985;
wire   [15:0] sub_ln703_209_fu_2157_p2;
reg   [15:0] sub_ln703_209_reg_10990;
wire   [15:0] sub_ln703_210_fu_2162_p2;
reg   [15:0] sub_ln703_210_reg_10995;
wire   [15:0] sub_ln703_212_fu_2173_p2;
reg   [15:0] sub_ln703_212_reg_11000;
wire   [15:0] add_ln703_323_fu_2188_p2;
reg   [15:0] add_ln703_323_reg_11005;
wire   [15:0] sub_ln703_230_fu_2194_p2;
reg   [15:0] sub_ln703_230_reg_11010;
wire   [15:0] add_ln703_328_fu_2208_p2;
reg   [15:0] add_ln703_328_reg_11015;
wire   [15:0] sub_ln703_237_fu_2214_p2;
reg   [15:0] sub_ln703_237_reg_11020;
wire   [15:0] add_ln703_333_fu_2224_p2;
reg   [15:0] add_ln703_333_reg_11025;
wire   [15:0] add_ln703_341_fu_2230_p2;
reg   [15:0] add_ln703_341_reg_11030;
wire   [15:0] add_ln703_369_fu_2234_p2;
reg   [15:0] add_ln703_369_reg_11037;
reg   [15:0] add_ln703_369_reg_11037_pp0_iter7_reg;
wire   [15:0] sub_ln703_234_fu_2395_p2;
reg   [15:0] sub_ln703_234_reg_11046;
wire   [15:0] sub_ln703_246_fu_2477_p2;
reg   [15:0] sub_ln703_246_reg_11051;
wire   [15:0] sub_ln703_249_fu_2496_p2;
reg   [15:0] sub_ln703_249_reg_11056;
wire   [15:0] sub_ln703_250_fu_2501_p2;
reg   [15:0] sub_ln703_250_reg_11061;
wire   [15:0] sub_ln703_251_fu_2506_p2;
reg   [15:0] sub_ln703_251_reg_11066;
wire   [15:0] add_ln703_342_fu_2520_p2;
reg   [15:0] add_ln703_342_reg_11071;
wire   [15:0] sub_ln703_254_fu_2525_p2;
reg   [15:0] sub_ln703_254_reg_11076;
wire   [15:0] sub_ln703_256_fu_2534_p2;
reg   [15:0] sub_ln703_256_reg_11081;
wire   [15:0] sub_ln703_257_fu_2539_p2;
reg   [15:0] sub_ln703_257_reg_11086;
wire   [15:0] sub_ln703_261_fu_2569_p2;
reg   [15:0] sub_ln703_261_reg_11091;
wire   [15:0] sub_ln703_262_fu_2574_p2;
reg   [15:0] sub_ln703_262_reg_11096;
wire   [15:0] sub_ln703_263_fu_2579_p2;
reg   [15:0] sub_ln703_263_reg_11101;
wire   [15:0] add_ln703_346_fu_2589_p2;
reg   [15:0] add_ln703_346_reg_11106;
wire   [15:0] add_ln703_350_fu_2602_p2;
reg   [15:0] add_ln703_350_reg_11111;
wire   [15:0] sub_ln703_265_fu_2613_p2;
reg   [15:0] sub_ln703_265_reg_11116;
wire   [15:0] sub_ln703_270_fu_2628_p2;
reg   [15:0] sub_ln703_270_reg_11121;
wire   [15:0] add_ln703_352_fu_2633_p2;
reg   [15:0] add_ln703_352_reg_11126;
wire   [15:0] add_ln703_354_fu_2638_p2;
reg   [15:0] add_ln703_354_reg_11131;
wire   [15:0] sub_ln703_272_fu_2647_p2;
reg   [15:0] sub_ln703_272_reg_11138;
wire   [15:0] sub_ln703_274_fu_2652_p2;
reg   [15:0] sub_ln703_274_reg_11143;
wire   [15:0] add_ln703_356_fu_2657_p2;
reg   [15:0] add_ln703_356_reg_11148;
wire   [15:0] sub_ln703_275_fu_2662_p2;
reg   [15:0] sub_ln703_275_reg_11153;
wire   [15:0] add_ln703_360_fu_2677_p2;
reg   [15:0] add_ln703_360_reg_11158;
wire   [15:0] sub_ln703_281_fu_2688_p2;
reg   [15:0] sub_ln703_281_reg_11163;
wire   [15:0] sub_ln703_284_fu_2698_p2;
reg   [15:0] sub_ln703_284_reg_11168;
wire   [15:0] sub_ln703_289_fu_2703_p2;
reg   [15:0] sub_ln703_289_reg_11173;
wire   [15:0] sub_ln703_293_fu_2708_p2;
reg   [15:0] sub_ln703_293_reg_11178;
wire   [15:0] sub_ln703_296_fu_2713_p2;
reg   [15:0] sub_ln703_296_reg_11183;
wire   [15:0] sub_ln703_301_fu_2718_p2;
reg   [15:0] sub_ln703_301_reg_11188;
wire   [15:0] add_ln703_371_fu_2732_p2;
reg   [15:0] add_ln703_371_reg_11193;
wire   [15:0] add_ln703_375_fu_2738_p2;
reg   [15:0] add_ln703_375_reg_11198;
wire   [15:0] add_ln703_384_fu_2743_p2;
reg   [15:0] add_ln703_384_reg_11203;
wire   [15:0] add_ln703_400_fu_2752_p2;
reg   [15:0] add_ln703_400_reg_11210;
wire   [15:0] add_ln703_402_fu_2758_p2;
reg   [15:0] add_ln703_402_reg_11215;
reg   [15:0] add_ln703_402_reg_11215_pp0_iter8_reg;
wire   [15:0] add_ln703_424_fu_2762_p2;
reg   [15:0] add_ln703_424_reg_11225;
wire   [15:0] add_ln703_439_fu_2766_p2;
reg   [15:0] add_ln703_439_reg_11233;
reg   [15:0] add_ln703_439_reg_11233_pp0_iter8_reg;
wire   [15:0] add_ln703_525_fu_2774_p2;
reg   [15:0] add_ln703_525_reg_11243;
reg   [15:0] add_ln703_525_reg_11243_pp0_iter8_reg;
reg   [15:0] add_ln703_525_reg_11243_pp0_iter9_reg;
wire   [15:0] add_ln703_534_fu_2779_p2;
reg   [15:0] add_ln703_534_reg_11248;
reg   [15:0] add_ln703_534_reg_11248_pp0_iter8_reg;
reg   [15:0] add_ln703_534_reg_11248_pp0_iter9_reg;
wire   [15:0] sub_ln703_313_fu_2998_p2;
reg   [15:0] sub_ln703_313_reg_11257;
wire   [15:0] add_ln703_386_fu_3015_p2;
reg   [15:0] add_ln703_386_reg_11262;
wire   [15:0] sub_ln703_315_fu_3021_p2;
reg   [15:0] sub_ln703_315_reg_11267;
wire   [15:0] add_ln703_390_fu_3050_p2;
reg   [15:0] add_ln703_390_reg_11272;
wire   [15:0] sub_ln703_326_fu_3101_p2;
reg   [15:0] sub_ln703_326_reg_11277;
wire   [15:0] sub_ln703_328_fu_3111_p2;
reg   [15:0] sub_ln703_328_reg_11282;
wire   [15:0] add_ln703_410_fu_3149_p2;
reg   [15:0] add_ln703_410_reg_11287;
wire   [15:0] sub_ln703_333_fu_3155_p2;
reg   [15:0] sub_ln703_333_reg_11292;
wire   [15:0] add_ln703_416_fu_3170_p2;
reg   [15:0] add_ln703_416_reg_11297;
wire   [15:0] sub_ln703_334_fu_3175_p2;
reg   [15:0] sub_ln703_334_reg_11302;
wire   [15:0] sub_ln703_336_fu_3180_p2;
reg   [15:0] sub_ln703_336_reg_11307;
wire   [15:0] add_ln703_417_fu_3185_p2;
reg   [15:0] add_ln703_417_reg_11312;
wire   [15:0] sub_ln703_339_fu_3200_p2;
reg   [15:0] sub_ln703_339_reg_11317;
wire   [15:0] sub_ln703_340_fu_3205_p2;
reg   [15:0] sub_ln703_340_reg_11322;
wire   [15:0] sub_ln703_342_fu_3215_p2;
reg   [15:0] sub_ln703_342_reg_11327;
wire   [15:0] sub_ln703_344_fu_3220_p2;
reg   [15:0] sub_ln703_344_reg_11332;
wire   [15:0] sub_ln703_345_fu_3234_p2;
reg   [15:0] sub_ln703_345_reg_11337;
wire   [15:0] sub_ln703_350_fu_3244_p2;
reg   [15:0] sub_ln703_350_reg_11342;
wire   [15:0] add_ln703_426_fu_3258_p2;
reg   [15:0] add_ln703_426_reg_11347;
wire   [15:0] sub_ln703_353_fu_3269_p2;
reg   [15:0] sub_ln703_353_reg_11352;
wire   [15:0] add_ln703_431_fu_3274_p2;
reg   [15:0] add_ln703_431_reg_11357;
wire   [15:0] add_ln703_435_fu_3284_p2;
reg   [15:0] add_ln703_435_reg_11362;
wire   [15:0] sub_ln703_356_fu_3290_p2;
reg   [15:0] sub_ln703_356_reg_11367;
wire   [15:0] sub_ln703_358_fu_3300_p2;
reg   [15:0] sub_ln703_358_reg_11372;
wire   [15:0] sub_ln703_362_fu_3305_p2;
reg   [15:0] sub_ln703_362_reg_11377;
wire   [15:0] add_ln703_438_fu_3310_p2;
reg   [15:0] add_ln703_438_reg_11382;
wire   [15:0] add_ln703_445_fu_3315_p2;
reg   [15:0] add_ln703_445_reg_11387;
wire   [15:0] add_ln703_447_fu_3320_p2;
reg   [15:0] add_ln703_447_reg_11392;
wire   [15:0] sub_ln703_371_fu_3324_p2;
reg   [15:0] sub_ln703_371_reg_11397;
wire   [15:0] add_ln703_451_fu_3329_p2;
reg   [15:0] add_ln703_451_reg_11402;
wire   [15:0] add_ln703_466_fu_3333_p2;
reg   [15:0] add_ln703_466_reg_11410;
wire   [15:0] add_ln703_471_fu_3337_p2;
reg   [15:0] add_ln703_471_reg_11418;
wire   [15:0] add_ln703_484_fu_3342_p2;
reg   [15:0] add_ln703_484_reg_11423;
wire   [15:0] add_ln703_490_fu_3347_p2;
reg   [15:0] add_ln703_490_reg_11428;
wire   [15:0] add_ln703_498_fu_3351_p2;
reg   [15:0] add_ln703_498_reg_11436;
wire   [15:0] add_ln703_507_fu_3356_p2;
reg   [15:0] add_ln703_507_reg_11441;
reg   [15:0] add_ln703_507_reg_11441_pp0_iter9_reg;
wire   [15:0] add_ln703_528_fu_3360_p2;
reg   [15:0] add_ln703_528_reg_11452;
reg   [15:0] add_ln703_528_reg_11452_pp0_iter9_reg;
wire   [15:0] add_ln703_535_fu_3364_p2;
reg   [15:0] add_ln703_535_reg_11457;
wire   [15:0] add_ln703_568_fu_3368_p2;
reg   [15:0] add_ln703_568_reg_11464;
reg   [15:0] add_ln703_568_reg_11464_pp0_iter9_reg;
wire   [15:0] sub_ln703_384_fu_3645_p2;
reg   [15:0] sub_ln703_384_reg_11474;
wire   [15:0] add_ln703_469_fu_3655_p2;
reg   [15:0] add_ln703_469_reg_11479;
wire   [15:0] sub_ln703_386_fu_3660_p2;
reg   [15:0] sub_ln703_386_reg_11484;
wire   [15:0] sub_ln703_387_fu_3665_p2;
reg   [15:0] sub_ln703_387_reg_11489;
wire   [15:0] add_ln703_476_fu_3685_p2;
reg   [15:0] add_ln703_476_reg_11494;
wire   [15:0] sub_ln703_390_fu_3690_p2;
reg   [15:0] sub_ln703_390_reg_11499;
wire   [15:0] sub_ln703_393_fu_3705_p2;
reg   [15:0] sub_ln703_393_reg_11504;
wire   [15:0] sub_ln703_394_fu_3710_p2;
reg   [15:0] sub_ln703_394_reg_11509;
wire   [15:0] sub_ln703_395_fu_3720_p2;
reg   [15:0] sub_ln703_395_reg_11514;
wire   [15:0] add_ln703_478_fu_3730_p2;
reg   [15:0] add_ln703_478_reg_11519;
wire   [15:0] sub_ln703_399_fu_3761_p2;
reg   [15:0] sub_ln703_399_reg_11524;
wire   [15:0] sub_ln703_401_fu_3781_p2;
reg   [15:0] sub_ln703_401_reg_11529;
wire   [15:0] sub_ln703_402_fu_3786_p2;
reg   [15:0] sub_ln703_402_reg_11534;
wire   [15:0] sub_ln703_403_fu_3791_p2;
reg   [15:0] sub_ln703_403_reg_11539;
wire   [15:0] add_ln703_496_fu_3806_p2;
reg   [15:0] add_ln703_496_reg_11544;
wire   [15:0] add_ln703_497_fu_3811_p2;
reg   [15:0] add_ln703_497_reg_11549;
wire   [15:0] sub_ln703_405_fu_3816_p2;
reg   [15:0] sub_ln703_405_reg_11554;
wire   [15:0] add_ln703_506_fu_3839_p2;
reg   [15:0] add_ln703_506_reg_11559;
wire   [15:0] sub_ln703_408_fu_3845_p2;
reg   [15:0] sub_ln703_408_reg_11564;
wire   [15:0] sub_ln703_411_fu_3850_p2;
reg   [15:0] sub_ln703_411_reg_11569;
wire   [15:0] sub_ln703_412_fu_3855_p2;
reg   [15:0] sub_ln703_412_reg_11574;
wire   [15:0] sub_ln703_414_fu_3860_p2;
reg   [15:0] sub_ln703_414_reg_11579;
wire   [15:0] sub_ln703_416_fu_3865_p2;
reg   [15:0] sub_ln703_416_reg_11584;
wire   [15:0] add_ln703_512_fu_3878_p2;
reg   [15:0] add_ln703_512_reg_11589;
wire   [15:0] sub_ln703_419_fu_3884_p2;
reg   [15:0] sub_ln703_419_reg_11594;
wire   [15:0] add_ln703_515_fu_3889_p2;
reg   [15:0] add_ln703_515_reg_11599;
wire   [15:0] add_ln703_517_fu_3894_p2;
reg   [15:0] add_ln703_517_reg_11604;
wire   [15:0] add_ln703_537_fu_3912_p2;
reg   [15:0] add_ln703_537_reg_11609;
wire   [15:0] add_ln703_545_fu_3923_p2;
reg   [15:0] add_ln703_545_reg_11614;
wire   [15:0] add_ln703_556_fu_3933_p2;
reg   [15:0] add_ln703_556_reg_11619;
wire   [15:0] sub_ln703_440_fu_3938_p2;
reg   [15:0] sub_ln703_440_reg_11624;
wire   [15:0] add_ln703_560_fu_3943_p2;
reg   [15:0] add_ln703_560_reg_11629;
wire   [15:0] add_ln703_566_fu_3952_p2;
reg   [15:0] add_ln703_566_reg_11635;
wire   [15:0] add_ln703_569_fu_3957_p2;
reg   [15:0] add_ln703_569_reg_11640;
wire   [15:0] add_ln703_588_fu_3961_p2;
reg   [15:0] add_ln703_588_reg_11646;
wire   [15:0] add_ln703_600_fu_3965_p2;
reg   [15:0] add_ln703_600_reg_11652;
reg   [15:0] add_ln703_600_reg_11652_pp0_iter10_reg;
wire   [15:0] add_ln703_621_fu_3969_p2;
reg   [15:0] add_ln703_621_reg_11662;
reg   [15:0] add_ln703_621_reg_11662_pp0_iter10_reg;
wire   [15:0] sub_ln703_448_fu_4206_p2;
reg   [15:0] sub_ln703_448_reg_11673;
wire   [15:0] sub_ln703_452_fu_4231_p2;
reg   [15:0] sub_ln703_452_reg_11678;
wire   [15:0] sub_ln703_453_fu_4236_p2;
reg   [15:0] sub_ln703_453_reg_11683;
wire   [15:0] sub_ln703_458_fu_4270_p2;
reg   [15:0] sub_ln703_458_reg_11688;
wire   [15:0] sub_ln703_461_fu_4303_p2;
reg   [15:0] sub_ln703_461_reg_11693;
wire   [15:0] add_ln703_572_fu_4308_p2;
reg   [15:0] add_ln703_572_reg_11698;
wire   [15:0] sub_ln703_462_fu_4313_p2;
reg   [15:0] sub_ln703_462_reg_11703;
wire   [15:0] add_ln703_573_fu_4323_p2;
reg   [15:0] add_ln703_573_reg_11708;
wire   [15:0] sub_ln703_467_fu_4333_p2;
reg   [15:0] sub_ln703_467_reg_11713;
wire   [15:0] sub_ln703_468_fu_4353_p2;
reg   [15:0] sub_ln703_468_reg_11718;
wire   [15:0] add_ln703_581_fu_4358_p2;
reg   [15:0] add_ln703_581_reg_11723;
wire   [15:0] add_ln703_583_fu_4363_p2;
reg   [15:0] add_ln703_583_reg_11728;
wire   [15:0] sub_ln703_469_fu_4368_p2;
reg   [15:0] sub_ln703_469_reg_11733;
wire   [15:0] sub_ln703_470_fu_4373_p2;
reg   [15:0] sub_ln703_470_reg_11738;
wire   [15:0] add_ln703_586_fu_4398_p2;
reg   [15:0] add_ln703_586_reg_11743;
wire   [15:0] add_ln703_590_fu_4412_p2;
reg   [15:0] add_ln703_590_reg_11748;
wire   [15:0] sub_ln703_475_fu_4418_p2;
reg   [15:0] sub_ln703_475_reg_11753;
wire   [15:0] add_ln703_591_fu_4423_p2;
reg   [15:0] add_ln703_591_reg_11758;
wire   [15:0] add_ln703_592_fu_4428_p2;
reg   [15:0] add_ln703_592_reg_11763;
wire   [15:0] add_ln703_598_fu_4441_p2;
reg   [15:0] add_ln703_598_reg_11768;
wire   [15:0] sub_ln703_482_fu_4447_p2;
reg   [15:0] sub_ln703_482_reg_11773;
wire   [15:0] sub_ln703_483_fu_4452_p2;
reg   [15:0] sub_ln703_483_reg_11778;
wire   [15:0] sub_ln703_488_fu_4457_p2;
reg   [15:0] sub_ln703_488_reg_11783;
wire   [15:0] sub_ln703_490_fu_4462_p2;
reg   [15:0] sub_ln703_490_reg_11788;
wire   [15:0] sub_ln703_491_fu_4467_p2;
reg   [15:0] sub_ln703_491_reg_11793;
wire   [15:0] add_ln703_599_fu_4477_p2;
reg   [15:0] add_ln703_599_reg_11798;
wire   [15:0] add_ln703_609_fu_4501_p2;
reg   [15:0] add_ln703_609_reg_11803;
wire   [15:0] add_ln703_616_fu_4511_p2;
reg   [15:0] add_ln703_616_reg_11808;
wire   [15:0] sub_ln703_503_fu_4516_p2;
reg   [15:0] sub_ln703_503_reg_11813;
wire   [15:0] sub_ln703_505_fu_4521_p2;
reg   [15:0] sub_ln703_505_reg_11818;
wire   [15:0] add_ln703_633_fu_4531_p2;
reg   [15:0] add_ln703_633_reg_11823;
wire   [15:0] add_ln703_634_fu_4535_p2;
reg   [15:0] add_ln703_634_reg_11828;
wire   [15:0] add_ln703_639_fu_4541_p2;
reg   [15:0] add_ln703_639_reg_11833;
wire   [15:0] add_ln703_646_fu_4546_p2;
reg   [15:0] add_ln703_646_reg_11838;
wire   [15:0] add_ln703_650_fu_4550_p2;
reg   [15:0] add_ln703_650_reg_11844;
reg   [15:0] add_ln703_650_reg_11844_pp0_iter11_reg;
wire   [15:0] add_ln703_667_fu_4554_p2;
reg   [15:0] add_ln703_667_reg_11853;
wire   [15:0] sub_ln703_526_fu_4860_p2;
reg   [15:0] sub_ln703_526_reg_11864;
wire   [15:0] sub_ln703_527_fu_4865_p2;
reg   [15:0] sub_ln703_527_reg_11869;
wire   [15:0] add_ln703_647_fu_4870_p2;
reg   [15:0] add_ln703_647_reg_11874;
wire   [15:0] sub_ln703_529_fu_4880_p2;
reg   [15:0] sub_ln703_529_reg_11879;
wire   [15:0] sub_ln703_532_fu_4894_p2;
reg   [15:0] sub_ln703_532_reg_11884;
wire   [15:0] add_ln703_648_fu_4899_p2;
reg   [15:0] add_ln703_648_reg_11889;
wire   [15:0] sub_ln703_533_fu_4904_p2;
reg   [15:0] sub_ln703_533_reg_11894;
wire   [15:0] sub_ln703_535_fu_4919_p2;
reg   [15:0] sub_ln703_535_reg_11899;
wire   [15:0] sub_ln703_538_fu_4934_p2;
reg   [15:0] sub_ln703_538_reg_11904;
wire   [15:0] sub_ln703_539_fu_4939_p2;
reg   [15:0] sub_ln703_539_reg_11909;
wire   [15:0] sub_ln703_540_fu_4944_p2;
reg   [15:0] sub_ln703_540_reg_11914;
wire   [15:0] sub_ln703_541_fu_4949_p2;
reg   [15:0] sub_ln703_541_reg_11919;
wire   [15:0] sub_ln703_542_fu_4954_p2;
reg   [15:0] sub_ln703_542_reg_11924;
wire   [15:0] add_ln703_651_fu_4959_p2;
reg   [15:0] add_ln703_651_reg_11929;
wire   [15:0] sub_ln703_544_fu_4984_p2;
reg   [15:0] sub_ln703_544_reg_11934;
wire   [15:0] add_ln703_660_fu_4994_p2;
reg   [15:0] add_ln703_660_reg_11939;
wire   [15:0] add_ln703_661_fu_4999_p2;
reg   [15:0] add_ln703_661_reg_11944;
wire   [15:0] sub_ln703_551_fu_5004_p2;
reg   [15:0] sub_ln703_551_reg_11949;
wire   [15:0] add_ln703_666_fu_5013_p2;
reg   [15:0] add_ln703_666_reg_11954;
wire   [15:0] add_ln703_668_fu_5019_p2;
reg   [15:0] add_ln703_668_reg_11959;
wire   [15:0] sub_ln703_556_fu_5024_p2;
reg   [15:0] sub_ln703_556_reg_11964;
wire   [15:0] sub_ln703_557_fu_5029_p2;
reg   [15:0] sub_ln703_557_reg_11969;
wire   [15:0] sub_ln703_558_fu_5034_p2;
reg   [15:0] sub_ln703_558_reg_11974;
wire   [15:0] add_ln703_676_fu_5052_p2;
reg   [15:0] add_ln703_676_reg_11979;
wire   [15:0] add_ln703_682_fu_5066_p2;
reg   [15:0] add_ln703_682_reg_11984;
wire   [15:0] add_ln703_685_fu_5077_p2;
reg   [15:0] add_ln703_685_reg_11989;
wire   [15:0] add_ln703_691_fu_5092_p2;
reg   [15:0] add_ln703_691_reg_11994;
wire   [15:0] add_ln703_697_fu_5096_p2;
reg   [15:0] add_ln703_697_reg_12002;
wire   [15:0] sub_ln703_573_fu_5101_p2;
reg   [15:0] sub_ln703_573_reg_12007;
wire   [15:0] sub_ln703_582_fu_5106_p2;
reg   [15:0] sub_ln703_582_reg_12012;
wire   [15:0] sub_ln703_583_fu_5111_p2;
reg   [15:0] sub_ln703_583_reg_12017;
wire   [15:0] add_ln703_703_fu_5116_p2;
reg   [15:0] add_ln703_703_reg_12022;
wire   [15:0] add_ln703_706_fu_5120_p2;
reg   [15:0] add_ln703_706_reg_12031;
wire   [15:0] add_ln703_722_fu_5125_p2;
reg   [15:0] add_ln703_722_reg_12036;
wire   [15:0] add_ln703_726_fu_5130_p2;
reg   [15:0] add_ln703_726_reg_12041;
wire   [15:0] add_ln703_737_fu_5134_p2;
reg   [15:0] add_ln703_737_reg_12047;
wire   [15:0] add_ln703_704_fu_5336_p2;
reg   [15:0] add_ln703_704_reg_12056;
wire   [15:0] sub_ln703_586_fu_5351_p2;
reg   [15:0] sub_ln703_586_reg_12061;
wire   [15:0] sub_ln703_589_fu_5375_p2;
reg   [15:0] sub_ln703_589_reg_12066;
wire   [15:0] sub_ln703_593_fu_5410_p2;
reg   [15:0] sub_ln703_593_reg_12071;
wire   [15:0] sub_ln703_594_fu_5415_p2;
reg   [15:0] sub_ln703_594_reg_12076;
wire   [15:0] sub_ln703_595_fu_5420_p2;
reg   [15:0] sub_ln703_595_reg_12081;
wire   [15:0] add_ln703_719_fu_5439_p2;
reg   [15:0] add_ln703_719_reg_12086;
wire   [15:0] sub_ln703_598_fu_5454_p2;
reg   [15:0] sub_ln703_598_reg_12091;
wire   [15:0] add_ln703_728_fu_5485_p2;
reg   [15:0] add_ln703_728_reg_12096;
wire   [15:0] sub_ln703_603_fu_5491_p2;
reg   [15:0] sub_ln703_603_reg_12101;
wire   [15:0] sub_ln703_604_fu_5496_p2;
reg   [15:0] sub_ln703_604_reg_12106;
wire   [15:0] sub_ln703_605_fu_5501_p2;
reg   [15:0] sub_ln703_605_reg_12111;
wire   [15:0] sub_ln703_608_fu_5511_p2;
reg   [15:0] sub_ln703_608_reg_12116;
wire   [15:0] sub_ln703_609_fu_5516_p2;
reg   [15:0] sub_ln703_609_reg_12121;
wire   [15:0] sub_ln703_610_fu_5521_p2;
reg   [15:0] sub_ln703_610_reg_12126;
wire   [15:0] sub_ln703_612_fu_5526_p2;
reg   [15:0] sub_ln703_612_reg_12131;
wire   [15:0] sub_ln703_613_fu_5531_p2;
reg   [15:0] sub_ln703_613_reg_12136;
wire   [15:0] sub_ln703_614_fu_5536_p2;
reg   [15:0] sub_ln703_614_reg_12141;
wire   [15:0] add_ln703_733_fu_5551_p2;
reg   [15:0] add_ln703_733_reg_12146;
wire   [15:0] add_ln703_734_fu_5556_p2;
reg   [15:0] add_ln703_734_reg_12151;
wire   [15:0] sub_ln703_618_fu_5566_p2;
reg   [15:0] sub_ln703_618_reg_12156;
wire   [15:0] add_ln703_735_fu_5571_p2;
reg   [15:0] add_ln703_735_reg_12161;
wire   [15:0] sub_ln703_624_fu_5596_p2;
reg   [15:0] sub_ln703_624_reg_12166;
wire   [15:0] sub_ln703_630_fu_5627_p2;
reg   [15:0] sub_ln703_630_reg_12171;
wire   [15:0] sub_ln703_631_fu_5632_p2;
reg   [15:0] sub_ln703_631_reg_12176;
wire   [15:0] sub_ln703_634_fu_5637_p2;
reg   [15:0] sub_ln703_634_reg_12181;
wire   [15:0] sub_ln703_637_fu_5642_p2;
reg   [15:0] sub_ln703_637_reg_12186;
wire   [15:0] sub_ln703_638_fu_5647_p2;
reg   [15:0] sub_ln703_638_reg_12191;
wire   [15:0] add_ln703_755_fu_5652_p2;
reg   [15:0] add_ln703_755_reg_12196;
wire   [15:0] sub_ln703_644_fu_5656_p2;
reg   [15:0] sub_ln703_644_reg_12204;
wire   [15:0] sub_ln703_648_fu_5661_p2;
reg   [15:0] sub_ln703_648_reg_12209;
wire   [15:0] sub_ln703_650_fu_5666_p2;
reg   [15:0] sub_ln703_650_reg_12214;
wire   [15:0] add_ln703_765_fu_5671_p2;
reg   [15:0] add_ln703_765_reg_12219;
wire   [15:0] add_ln703_778_fu_5675_p2;
reg   [15:0] add_ln703_778_reg_12227;
wire   [15:0] add_ln703_783_fu_5679_p2;
reg   [15:0] add_ln703_783_reg_12236;
wire   [15:0] add_ln703_816_fu_5684_p2;
reg   [15:0] add_ln703_816_reg_12241;
reg   [15:0] add_ln703_816_reg_12241_pp0_iter13_reg;
wire   [15:0] sub_ln703_662_fu_5918_p2;
reg   [15:0] sub_ln703_662_reg_12248;
wire   [15:0] sub_ln703_665_fu_5932_p2;
reg   [15:0] sub_ln703_665_reg_12253;
wire   [15:0] add_ln703_770_fu_5950_p2;
reg   [15:0] add_ln703_770_reg_12258;
wire   [15:0] sub_ln703_667_fu_5956_p2;
reg   [15:0] sub_ln703_667_reg_12263;
wire   [15:0] sub_ln703_669_fu_5975_p2;
reg   [15:0] sub_ln703_669_reg_12268;
wire   [15:0] add_ln703_779_fu_6024_p2;
reg   [15:0] add_ln703_779_reg_12273;
wire   [15:0] sub_ln703_676_fu_6033_p2;
reg   [15:0] sub_ln703_676_reg_12278;
wire   [15:0] sub_ln703_678_fu_6052_p2;
reg   [15:0] sub_ln703_678_reg_12283;
wire   [15:0] sub_ln703_679_fu_6057_p2;
reg   [15:0] sub_ln703_679_reg_12288;
wire   [15:0] sub_ln703_680_fu_6062_p2;
reg   [15:0] sub_ln703_680_reg_12293;
wire   [15:0] sub_ln703_682_fu_6067_p2;
reg   [15:0] sub_ln703_682_reg_12298;
wire   [15:0] sub_ln703_684_fu_6072_p2;
reg   [15:0] sub_ln703_684_reg_12303;
wire   [15:0] sub_ln703_686_fu_6077_p2;
reg   [15:0] sub_ln703_686_reg_12308;
wire   [15:0] sub_ln703_687_fu_6086_p2;
reg   [15:0] sub_ln703_687_reg_12313;
wire   [15:0] sub_ln703_688_fu_6091_p2;
reg   [15:0] sub_ln703_688_reg_12318;
wire   [15:0] sub_ln703_690_fu_6101_p2;
reg   [15:0] sub_ln703_690_reg_12323;
wire   [15:0] sub_ln703_691_fu_6106_p2;
reg   [15:0] sub_ln703_691_reg_12328;
wire   [15:0] sub_ln703_692_fu_6111_p2;
reg   [15:0] sub_ln703_692_reg_12333;
wire   [15:0] sub_ln703_693_fu_6116_p2;
reg   [15:0] sub_ln703_693_reg_12338;
wire   [15:0] sub_ln703_694_fu_6126_p2;
reg   [15:0] sub_ln703_694_reg_12343;
wire   [15:0] add_ln703_791_fu_6131_p2;
reg   [15:0] add_ln703_791_reg_12348;
wire   [15:0] sub_ln703_696_fu_6136_p2;
reg   [15:0] sub_ln703_696_reg_12353;
wire   [15:0] sub_ln703_697_fu_6141_p2;
reg   [15:0] sub_ln703_697_reg_12358;
wire   [15:0] add_ln703_792_fu_6146_p2;
reg   [15:0] add_ln703_792_reg_12363;
wire   [15:0] add_ln703_796_fu_6160_p2;
reg   [15:0] add_ln703_796_reg_12368;
wire   [15:0] add_ln703_798_fu_6166_p2;
reg   [15:0] add_ln703_798_reg_12373;
wire   [15:0] sub_ln703_700_fu_6172_p2;
reg   [15:0] sub_ln703_700_reg_12378;
wire   [15:0] sub_ln703_704_fu_6177_p2;
reg   [15:0] sub_ln703_704_reg_12383;
wire   [15:0] sub_ln703_707_fu_6182_p2;
reg   [15:0] sub_ln703_707_reg_12388;
wire   [15:0] add_ln703_801_fu_6187_p2;
reg   [15:0] add_ln703_801_reg_12393;
wire   [15:0] add_ln703_802_fu_6192_p2;
reg   [15:0] add_ln703_802_reg_12398;
wire   [15:0] add_ln703_818_fu_6205_p2;
reg   [15:0] add_ln703_818_reg_12409;
reg   [15:0] add_ln703_818_reg_12409_pp0_iter14_reg;
wire   [15:0] add_ln703_821_fu_6216_p2;
reg   [15:0] add_ln703_821_reg_12414;
wire   [15:0] add_ln703_826_fu_6222_p2;
reg   [15:0] add_ln703_826_reg_12419;
wire   [15:0] add_ln703_836_fu_6226_p2;
reg   [15:0] add_ln703_836_reg_12428;
wire   [15:0] add_ln703_849_fu_6230_p2;
reg   [15:0] add_ln703_849_reg_12434;
reg   [15:0] add_ln703_849_reg_12434_pp0_iter14_reg;
wire   [15:0] add_ln703_867_fu_6234_p2;
reg   [15:0] add_ln703_867_reg_12444;
reg   [15:0] add_ln703_867_reg_12444_pp0_iter14_reg;
wire   [15:0] sub_ln703_724_fu_6432_p2;
reg   [15:0] sub_ln703_724_reg_12450;
wire   [15:0] add_ln703_819_fu_6447_p2;
reg   [15:0] add_ln703_819_reg_12455;
wire   [15:0] sub_ln703_727_fu_6452_p2;
reg   [15:0] sub_ln703_727_reg_12460;
wire   [15:0] sub_ln703_728_fu_6457_p2;
reg   [15:0] sub_ln703_728_reg_12465;
wire   [15:0] sub_ln703_733_fu_6487_p2;
reg   [15:0] sub_ln703_733_reg_12470;
wire   [15:0] sub_ln703_736_fu_6502_p2;
reg   [15:0] sub_ln703_736_reg_12475;
wire   [15:0] add_ln703_825_fu_6526_p2;
reg   [15:0] add_ln703_825_reg_12480;
wire   [15:0] add_ln703_827_fu_6531_p2;
reg   [15:0] add_ln703_827_reg_12485;
wire   [15:0] add_ln703_831_fu_6554_p2;
reg   [15:0] add_ln703_831_reg_12490;
wire   [15:0] add_ln703_833_fu_6573_p2;
reg   [15:0] add_ln703_833_reg_12495;
wire   [15:0] sub_ln703_746_fu_6579_p2;
reg   [15:0] sub_ln703_746_reg_12500;
wire   [15:0] add_ln703_834_fu_6594_p2;
reg   [15:0] add_ln703_834_reg_12505;
wire   [15:0] sub_ln703_749_fu_6599_p2;
reg   [15:0] sub_ln703_749_reg_12510;
wire   [15:0] sub_ln703_757_fu_6629_p2;
reg   [15:0] sub_ln703_757_reg_12515;
wire   [15:0] add_ln703_838_fu_6634_p2;
reg   [15:0] add_ln703_838_reg_12520;
wire   [15:0] sub_ln703_759_fu_6639_p2;
reg   [15:0] sub_ln703_759_reg_12525;
wire   [15:0] sub_ln703_761_fu_6644_p2;
reg   [15:0] sub_ln703_761_reg_12530;
wire   [15:0] add_ln703_840_fu_6649_p2;
reg   [15:0] add_ln703_840_reg_12535;
wire   [15:0] sub_ln703_763_fu_6654_p2;
reg   [15:0] sub_ln703_763_reg_12540;
wire   [15:0] sub_ln703_767_fu_6659_p2;
reg   [15:0] sub_ln703_767_reg_12545;
wire   [15:0] add_ln703_841_fu_6664_p2;
reg   [15:0] add_ln703_841_reg_12550;
wire   [15:0] sub_ln703_769_fu_6684_p2;
reg   [15:0] sub_ln703_769_reg_12555;
wire   [15:0] add_ln703_845_fu_6689_p2;
reg   [15:0] add_ln703_845_reg_12560;
wire   [15:0] add_ln703_851_fu_6702_p2;
reg   [15:0] add_ln703_851_reg_12565;
wire   [15:0] sub_ln703_770_fu_6708_p2;
reg   [15:0] sub_ln703_770_reg_12570;
wire   [15:0] add_ln703_858_fu_6733_p2;
reg   [15:0] add_ln703_858_reg_12575;
wire   [15:0] sub_ln703_781_fu_6739_p2;
reg   [15:0] sub_ln703_781_reg_12580;
wire   [15:0] add_ln703_868_fu_6755_p2;
reg   [15:0] add_ln703_868_reg_12585;
wire   [15:0] sub_ln703_787_fu_6759_p2;
reg   [15:0] sub_ln703_787_reg_12590;
wire   [15:0] sub_ln703_799_fu_6764_p2;
reg   [15:0] sub_ln703_799_reg_12595;
wire   [15:0] add_ln703_876_fu_6769_p2;
reg   [15:0] add_ln703_876_reg_12600;
wire   [15:0] add_ln703_877_fu_6774_p2;
reg   [15:0] add_ln703_877_reg_12605;
wire   [15:0] add_ln703_894_fu_6778_p2;
reg   [15:0] add_ln703_894_reg_12616;
reg   [15:0] add_ln703_894_reg_12616_pp0_iter15_reg;
wire   [15:0] add_ln703_905_fu_6782_p2;
reg   [15:0] add_ln703_905_reg_12625;
wire   [15:0] add_ln703_914_fu_6786_p2;
reg   [15:0] add_ln703_914_reg_12632;
wire   [15:0] add_ln703_920_fu_6791_p2;
reg   [15:0] add_ln703_920_reg_12637;
reg   [15:0] add_ln703_920_reg_12637_pp0_iter15_reg;
wire   [15:0] sub_ln703_797_fu_7030_p2;
reg   [15:0] sub_ln703_797_reg_12645;
wire   [15:0] add_ln703_872_fu_7050_p2;
reg   [15:0] add_ln703_872_reg_12650;
wire   [15:0] add_ln703_873_fu_7055_p2;
reg   [15:0] add_ln703_873_reg_12655;
wire   [15:0] sub_ln703_801_fu_7060_p2;
reg   [15:0] sub_ln703_801_reg_12660;
wire   [15:0] sub_ln703_802_fu_7065_p2;
reg   [15:0] sub_ln703_802_reg_12665;
wire   [15:0] sub_ln703_805_fu_7079_p2;
reg   [15:0] sub_ln703_805_reg_12670;
wire   [15:0] add_ln703_874_fu_7084_p2;
reg   [15:0] add_ln703_874_reg_12675;
wire   [15:0] add_ln703_875_fu_7094_p2;
reg   [15:0] add_ln703_875_reg_12680;
wire   [15:0] sub_ln703_807_fu_7099_p2;
reg   [15:0] sub_ln703_807_reg_12685;
wire   [15:0] add_ln703_882_fu_7121_p2;
reg   [15:0] add_ln703_882_reg_12690;
wire   [15:0] add_ln703_884_fu_7132_p2;
reg   [15:0] add_ln703_884_reg_12695;
wire   [15:0] sub_ln703_808_fu_7137_p2;
reg   [15:0] sub_ln703_808_reg_12700;
wire   [15:0] add_ln703_888_fu_7156_p2;
reg   [15:0] add_ln703_888_reg_12705;
wire   [15:0] add_ln703_892_fu_7175_p2;
reg   [15:0] add_ln703_892_reg_12710;
wire   [15:0] add_ln703_893_fu_7180_p2;
reg   [15:0] add_ln703_893_reg_12715;
wire   [15:0] add_ln703_895_fu_7185_p2;
reg   [15:0] add_ln703_895_reg_12720;
wire   [15:0] add_ln703_896_fu_7190_p2;
reg   [15:0] add_ln703_896_reg_12725;
wire   [15:0] add_ln703_898_fu_7195_p2;
reg   [15:0] add_ln703_898_reg_12730;
wire   [15:0] sub_ln703_814_fu_7200_p2;
reg   [15:0] sub_ln703_814_reg_12735;
wire   [15:0] sub_ln703_816_fu_7205_p2;
reg   [15:0] sub_ln703_816_reg_12740;
wire   [15:0] sub_ln703_818_fu_7210_p2;
reg   [15:0] sub_ln703_818_reg_12745;
wire   [15:0] sub_ln703_820_fu_7215_p2;
reg   [15:0] sub_ln703_820_reg_12750;
wire   [15:0] sub_ln703_821_fu_7220_p2;
reg   [15:0] sub_ln703_821_reg_12755;
wire   [15:0] sub_ln703_823_fu_7225_p2;
reg   [15:0] sub_ln703_823_reg_12760;
wire   [15:0] sub_ln703_824_fu_7230_p2;
reg   [15:0] sub_ln703_824_reg_12765;
wire   [15:0] sub_ln703_825_fu_7235_p2;
reg   [15:0] sub_ln703_825_reg_12770;
wire   [15:0] add_ln703_906_fu_7245_p2;
reg   [15:0] add_ln703_906_reg_12775;
wire   [15:0] add_ln703_917_fu_7273_p2;
reg   [15:0] add_ln703_917_reg_12780;
wire   [15:0] add_ln703_922_fu_7287_p2;
reg   [15:0] add_ln703_922_reg_12785;
wire   [15:0] sub_ln703_852_fu_7319_p2;
reg   [15:0] sub_ln703_852_reg_12790;
wire   [15:0] sub_ln703_862_fu_7324_p2;
reg   [15:0] sub_ln703_862_reg_12795;
wire   [15:0] sub_ln703_869_fu_7329_p2;
reg   [15:0] sub_ln703_869_reg_12800;
reg   [15:0] sub_ln703_869_reg_12800_pp0_iter16_reg;
wire   [15:0] add_ln703_946_fu_7334_p2;
reg   [15:0] add_ln703_946_reg_12805;
wire   [15:0] add_ln703_954_fu_7338_p2;
reg   [15:0] add_ln703_954_reg_12812;
wire   [15:0] add_ln703_985_fu_7342_p2;
reg   [15:0] add_ln703_985_reg_12819;
reg   [15:0] add_ln703_985_reg_12819_pp0_iter16_reg;
wire   [15:0] sub_ln703_857_fu_7600_p2;
reg   [15:0] sub_ln703_857_reg_12835;
wire   [15:0] sub_ln703_858_fu_7605_p2;
reg   [15:0] sub_ln703_858_reg_12840;
wire   [15:0] add_ln703_934_fu_7610_p2;
reg   [15:0] add_ln703_934_reg_12845;
wire   [15:0] sub_ln703_859_fu_7615_p2;
reg   [15:0] sub_ln703_859_reg_12850;
wire   [15:0] add_ln703_936_fu_7634_p2;
reg   [15:0] add_ln703_936_reg_12855;
wire   [15:0] sub_ln703_863_fu_7639_p2;
reg   [15:0] sub_ln703_863_reg_12860;
wire   [15:0] sub_ln703_865_fu_7649_p2;
reg   [15:0] sub_ln703_865_reg_12865;
wire   [15:0] sub_ln703_866_fu_7654_p2;
reg   [15:0] sub_ln703_866_reg_12870;
wire   [15:0] add_ln703_938_fu_7663_p2;
reg   [15:0] add_ln703_938_reg_12875;
wire   [15:0] sub_ln703_867_fu_7669_p2;
reg   [15:0] sub_ln703_867_reg_12880;
wire   [15:0] sub_ln703_868_fu_7674_p2;
reg   [15:0] sub_ln703_868_reg_12885;
wire   [15:0] add_ln703_939_fu_7679_p2;
reg   [15:0] add_ln703_939_reg_12890;
wire   [15:0] sub_ln703_870_fu_7685_p2;
reg   [15:0] sub_ln703_870_reg_12895;
wire   [15:0] sub_ln703_873_fu_7710_p2;
reg   [15:0] sub_ln703_873_reg_12900;
wire   [15:0] add_ln703_943_fu_7719_p2;
reg   [15:0] add_ln703_943_reg_12905;
wire   [15:0] sub_ln703_875_fu_7730_p2;
reg   [15:0] sub_ln703_875_reg_12910;
wire   [15:0] sub_ln703_879_fu_7735_p2;
reg   [15:0] sub_ln703_879_reg_12915;
wire   [15:0] sub_ln703_880_fu_7750_p2;
reg   [15:0] sub_ln703_880_reg_12920;
wire   [15:0] sub_ln703_881_fu_7755_p2;
reg   [15:0] sub_ln703_881_reg_12925;
wire   [15:0] add_ln703_948_fu_7760_p2;
reg   [15:0] add_ln703_948_reg_12930;
wire   [15:0] sub_ln703_892_fu_7780_p2;
reg   [15:0] sub_ln703_892_reg_12935;
wire   [15:0] sub_ln703_893_fu_7785_p2;
reg   [15:0] sub_ln703_893_reg_12940;
wire   [15:0] sub_ln703_894_fu_7790_p2;
reg   [15:0] sub_ln703_894_reg_12945;
wire   [15:0] sub_ln703_895_fu_7795_p2;
reg   [15:0] sub_ln703_895_reg_12950;
wire   [15:0] sub_ln703_898_fu_7805_p2;
reg   [15:0] sub_ln703_898_reg_12955;
wire   [15:0] sub_ln703_904_fu_7810_p2;
reg   [15:0] sub_ln703_904_reg_12960;
wire   [15:0] add_ln703_958_fu_7827_p2;
reg   [15:0] add_ln703_958_reg_12965;
wire   [15:0] sub_ln703_911_fu_7833_p2;
reg   [15:0] sub_ln703_911_reg_12970;
wire   [15:0] sub_ln703_917_fu_7838_p2;
reg   [15:0] sub_ln703_917_reg_12975;
wire   [15:0] sub_ln703_922_fu_7843_p2;
reg   [15:0] sub_ln703_922_reg_12980;
wire   [15:0] add_ln703_964_fu_7848_p2;
reg   [15:0] add_ln703_964_reg_12985;
wire   [15:0] acc_21_V_fu_7872_p2;
reg   [15:0] acc_21_V_reg_12991;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_5_fu_564_p2;
wire   [15:0] add_ln703_143_fu_585_p2;
wire   [15:0] add_ln703_142_fu_581_p2;
wire   [15:0] add_ln703_133_fu_603_p2;
wire   [15:0] sub_ln703_7_fu_607_p2;
wire   [15:0] sub_ln703_9_fu_611_p2;
wire   [15:0] add_ln703_136_fu_623_p2;
wire   [15:0] add_ln703_139_fu_636_p2;
wire   [15:0] sub_ln703_12_fu_627_p2;
wire   [15:0] sub_ln703_13_fu_689_p2;
wire   [15:0] sub_ln703_14_fu_693_p2;
wire   [15:0] add_ln703_137_fu_697_p2;
wire   [15:0] add_ln703_138_fu_701_p2;
wire   [15:0] sub_ln703_19_fu_705_p2;
wire   [15:0] sub_ln703_22_fu_713_p2;
wire   [15:0] sub_ln703_24_fu_717_p2;
wire   [15:0] sub_ln703_25_fu_722_p2;
wire   [15:0] sub_ln703_27_fu_732_p2;
wire   [15:0] add_ln703_145_fu_736_p2;
wire   [15:0] add_ln703_146_fu_741_p2;
wire   [15:0] add_ln703_147_fu_745_p2;
wire   [15:0] sub_ln703_29_fu_749_p2;
wire   [15:0] sub_ln703_30_fu_753_p2;
wire   [15:0] add_ln703_148_fu_757_p2;
wire   [15:0] sub_ln703_31_fu_761_p2;
wire   [15:0] sub_ln703_32_fu_765_p2;
wire   [15:0] sub_ln703_33_fu_769_p2;
wire   [15:0] add_ln703_155_fu_868_p2;
wire   [15:0] add_ln703_149_fu_773_p2;
wire   [15:0] sub_ln703_34_fu_778_p2;
wire   [15:0] add_ln703_150_fu_782_p2;
wire   [15:0] sub_ln703_35_fu_787_p2;
wire   [15:0] add_ln703_151_fu_791_p2;
wire   [15:0] sub_ln703_37_fu_800_p2;
wire   [15:0] add_ln703_152_fu_804_p2;
wire   [15:0] sub_ln703_26_fu_727_p2;
wire   [15:0] sub_ln703_41_fu_829_p2;
wire   [15:0] add_ln703_154_fu_843_p2;
wire   [15:0] sub_ln703_44_fu_848_p2;
wire   [15:0] sub_ln703_45_fu_853_p2;
wire   [15:0] add_ln703_156_fu_872_p2;
wire   [15:0] sub_ln703_48_fu_877_p2;
wire   [15:0] sub_ln703_49_fu_882_p2;
wire   [15:0] sub_ln703_21_fu_709_p2;
wire   [15:0] add_ln703_166_fu_962_p2;
wire   [15:0] sub_ln703_51_fu_897_p2;
wire   [15:0] sub_ln703_36_fu_795_p2;
wire   [15:0] add_ln703_160_fu_902_p2;
wire   [15:0] sub_ln703_60_fu_927_p2;
wire   [15:0] sub_ln703_61_fu_932_p2;
wire   [15:0] add_ln703_164_fu_937_p2;
wire   [15:0] add_ln703_180_fu_1011_p2;
wire   [15:0] add_ln703_178_fu_1007_p2;
wire   [15:0] sub_ln703_47_fu_863_p2;
wire   [15:0] add_ln703_165_fu_952_p2;
wire   [15:0] add_ln703_168_fu_967_p2;
wire   [15:0] sub_ln703_50_fu_887_p2;
wire   [15:0] add_ln703_187_fu_1041_p2;
wire   [15:0] add_ln703_189_fu_1045_p2;
wire   [15:0] sub_ln703_52_fu_907_p2;
wire   [15:0] sub_ln703_46_fu_858_p2;
wire   [15:0] sub_ln703_42_fu_833_p2;
wire   [15:0] sub_ln703_54_fu_1086_p2;
wire   [15:0] sub_ln703_55_fu_1090_p2;
wire   [15:0] sub_ln703_56_fu_1094_p2;
wire   [15:0] add_ln703_163_fu_1098_p2;
wire   [15:0] sub_ln703_57_fu_1102_p2;
wire   [15:0] sub_ln703_65_fu_1110_p2;
wire   [15:0] add_ln703_174_fu_1114_p2;
wire   [15:0] sub_ln703_67_fu_1119_p2;
wire   [15:0] add_ln703_175_fu_1123_p2;
wire   [15:0] add_ln703_176_fu_1128_p2;
wire   [15:0] sub_ln703_69_fu_1138_p2;
wire   [15:0] sub_ln703_59_fu_1106_p2;
wire   [15:0] add_ln703_184_fu_1143_p2;
wire   [15:0] sub_ln703_72_fu_1147_p2;
wire   [15:0] sub_ln703_74_fu_1151_p2;
wire   [15:0] sub_ln703_77_fu_1159_p2;
wire   [15:0] sub_ln703_78_fu_1164_p2;
wire   [15:0] sub_ln703_79_fu_1168_p2;
wire   [15:0] add_ln703_190_fu_1172_p2;
wire   [15:0] add_ln703_191_fu_1176_p2;
wire   [15:0] add_ln703_193_fu_1180_p2;
wire   [15:0] sub_ln703_80_fu_1184_p2;
wire   [15:0] add_ln703_194_fu_1189_p2;
wire   [15:0] sub_ln703_82_fu_1199_p2;
wire   [15:0] sub_ln703_68_fu_1133_p2;
wire   [15:0] add_ln703_195_fu_1204_p2;
wire   [15:0] add_ln703_197_fu_1209_p2;
wire   [15:0] add_ln703_199_fu_1213_p2;
wire   [15:0] sub_ln703_83_fu_1218_p2;
wire   [15:0] sub_ln703_84_fu_1222_p2;
wire   [15:0] add_ln703_200_fu_1226_p2;
wire   [15:0] add_ln703_214_fu_1349_p2;
wire   [15:0] sub_ln703_85_fu_1230_p2;
wire   [15:0] sub_ln703_87_fu_1238_p2;
wire   [15:0] add_ln703_201_fu_1243_p2;
wire   [15:0] sub_ln703_88_fu_1248_p2;
wire   [15:0] sub_ln703_89_fu_1252_p2;
wire   [15:0] sub_ln703_90_fu_1257_p2;
wire   [15:0] sub_ln703_91_fu_1261_p2;
wire   [15:0] add_ln703_217_fu_1393_p2;
wire   [15:0] sub_ln703_76_fu_1155_p2;
wire   [15:0] add_ln703_202_fu_1265_p2;
wire   [15:0] add_ln703_203_fu_1270_p2;
wire   [15:0] sub_ln703_93_fu_1275_p2;
wire   [15:0] sub_ln703_94_fu_1280_p2;
wire   [15:0] add_ln703_206_fu_1290_p2;
wire   [15:0] sub_ln703_97_fu_1304_p2;
wire   [15:0] sub_ln703_81_fu_1194_p2;
wire   [15:0] sub_ln703_99_fu_1324_p2;
wire   [15:0] add_ln703_211_fu_1339_p2;
wire   [15:0] sub_ln703_102_fu_1344_p2;
wire   [15:0] add_ln703_215_fu_1353_p2;
wire   [15:0] sub_ln703_103_fu_1363_p2;
wire   [15:0] sub_ln703_104_fu_1368_p2;
wire   [15:0] sub_ln703_105_fu_1373_p2;
wire   [15:0] add_ln703_219_fu_1397_p2;
wire   [15:0] add_ln703_221_fu_1402_p2;
wire   [15:0] sub_ln703_111_fu_1417_p2;
wire   [15:0] sub_ln703_112_fu_1422_p2;
wire   [15:0] sub_ln703_113_fu_1427_p2;
wire   [15:0] sub_ln703_119_fu_1442_p2;
wire   [15:0] add_ln703_237_fu_1516_p2;
wire   [15:0] sub_ln703_100_fu_1329_p2;
wire   [15:0] sub_ln703_101_fu_1334_p2;
wire   [15:0] add_ln703_225_fu_1452_p2;
wire   [15:0] sub_ln703_86_fu_1234_p2;
wire   [15:0] add_ln703_242_fu_1537_p2;
wire   [15:0] add_ln703_228_fu_1477_p2;
wire   [15:0] sub_ln703_126_fu_1487_p2;
wire   [15:0] add_ln703_232_fu_1492_p2;
wire   [15:0] sub_ln703_110_fu_1412_p2;
wire   [15:0] sub_ln703_95_fu_1285_p2;
wire   [15:0] add_ln703_248_fu_1569_p2;
wire   [15:0] sub_ln703_129_fu_1506_p2;
wire   [15:0] add_ln703_259_fu_1589_p2;
wire   [15:0] add_ln703_256_fu_1585_p2;
wire   [15:0] add_ln703_240_fu_1526_p2;
wire   [15:0] sub_ln703_120_fu_1447_p2;
wire   [15:0] add_ln703_244_fu_1542_p2;
wire   [15:0] add_ln703_222_fu_1626_p2;
wire   [15:0] sub_ln703_114_fu_1630_p2;
wire   [15:0] sub_ln703_118_fu_1642_p2;
wire   [15:0] sub_ln703_121_fu_1646_p2;
wire   [15:0] sub_ln703_124_fu_1650_p2;
wire   [15:0] add_ln703_229_fu_1654_p2;
wire   [15:0] add_ln703_230_fu_1658_p2;
wire   [15:0] sub_ln703_127_fu_1662_p2;
wire   [15:0] sub_ln703_130_fu_1666_p2;
wire   [15:0] add_ln703_234_fu_1671_p2;
wire   [15:0] add_ln703_235_fu_1676_p2;
wire   [15:0] sub_ln703_131_fu_1680_p2;
wire   [15:0] sub_ln703_117_fu_1638_p2;
wire   [15:0] add_ln703_241_fu_1693_p2;
wire   [15:0] sub_ln703_135_fu_1698_p2;
wire   [15:0] sub_ln703_136_fu_1702_p2;
wire   [15:0] sub_ln703_139_fu_1711_p2;
wire   [15:0] sub_ln703_140_fu_1716_p2;
wire   [15:0] add_ln703_245_fu_1721_p2;
wire   [15:0] sub_ln703_145_fu_1734_p2;
wire   [15:0] sub_ln703_148_fu_1743_p2;
wire   [15:0] sub_ln703_149_fu_1748_p2;
wire   [15:0] add_ln703_251_fu_1753_p2;
wire   [15:0] add_ln703_253_fu_1758_p2;
wire   [15:0] sub_ln703_132_fu_1684_p2;
wire   [15:0] sub_ln703_150_fu_1763_p2;
wire   [15:0] sub_ln703_151_fu_1767_p2;
wire   [15:0] add_ln703_263_fu_1771_p2;
wire   [15:0] sub_ln703_134_fu_1689_p2;
wire   [15:0] add_ln703_269_fu_1891_p2;
wire   [15:0] sub_ln703_156_fu_1785_p2;
wire   [15:0] sub_ln703_157_fu_1790_p2;
wire   [15:0] sub_ln703_138_fu_1706_p2;
wire   [15:0] sub_ln703_160_fu_1804_p2;
wire   [15:0] sub_ln703_161_fu_1809_p2;
wire   [15:0] sub_ln703_162_fu_1813_p2;
wire   [15:0] sub_ln703_143_fu_1725_p2;
wire   [15:0] sub_ln703_163_fu_1817_p2;
wire   [15:0] add_ln703_264_fu_1821_p2;
wire   [15:0] sub_ln703_164_fu_1826_p2;
wire   [15:0] sub_ln703_165_fu_1830_p2;
wire   [15:0] sub_ln703_168_fu_1844_p2;
wire   [15:0] sub_ln703_116_fu_1634_p2;
wire   [15:0] add_ln703_281_fu_1969_p2;
wire   [15:0] add_ln703_279_fu_1964_p2;
wire   [15:0] sub_ln703_169_fu_1849_p2;
wire   [15:0] add_ln703_266_fu_1854_p2;
wire   [15:0] sub_ln703_172_fu_1868_p2;
wire   [15:0] sub_ln703_173_fu_1873_p2;
wire   [15:0] sub_ln703_174_fu_1877_p2;
wire   [15:0] add_ln703_268_fu_1886_p2;
wire   [15:0] sub_ln703_153_fu_1775_p2;
wire   [15:0] add_ln703_271_fu_1895_p2;
wire   [15:0] sub_ln703_155_fu_1780_p2;
wire   [15:0] sub_ln703_178_fu_1909_p2;
wire   [15:0] add_ln703_273_fu_1914_p2;
wire   [15:0] sub_ln703_158_fu_1794_p2;
wire   [15:0] sub_ln703_179_fu_1919_p2;
wire   [15:0] add_ln703_274_fu_1924_p2;
wire   [15:0] sub_ln703_180_fu_1929_p2;
wire   [15:0] add_ln703_276_fu_1934_p2;
wire   [15:0] add_ln703_277_fu_1939_p2;
wire   [15:0] sub_ln703_144_fu_1730_p2;
wire   [15:0] add_ln703_291_fu_2064_p2;
wire   [15:0] sub_ln703_181_fu_1944_p2;
wire   [15:0] add_ln703_278_fu_1954_p2;
wire   [15:0] sub_ln703_147_fu_1738_p2;
wire   [15:0] sub_ln703_167_fu_1839_p2;
wire   [15:0] add_ln703_282_fu_1973_p2;
wire   [15:0] sub_ln703_171_fu_1864_p2;
wire   [15:0] sub_ln703_185_fu_1989_p2;
wire   [15:0] sub_ln703_188_fu_2004_p2;
wire   [15:0] sub_ln703_189_fu_2014_p2;
wire   [15:0] sub_ln703_176_fu_1900_p2;
wire   [15:0] add_ln703_287_fu_2019_p2;
wire   [15:0] sub_ln703_177_fu_1904_p2;
wire   [15:0] sub_ln703_190_fu_2024_p2;
wire   [15:0] sub_ln703_159_fu_1799_p2;
wire   [15:0] sub_ln703_192_fu_2044_p2;
wire   [15:0] sub_ln703_195_fu_2059_p2;
wire   [15:0] add_ln703_293_fu_2069_p2;
wire   [15:0] sub_ln703_182_fu_1949_p2;
wire   [15:0] sub_ln703_197_fu_2079_p2;
wire   [15:0] add_ln703_316_fu_2178_p2;
wire   [15:0] sub_ln703_187_fu_1999_p2;
wire   [15:0] sub_ln703_193_fu_2049_p2;
wire   [15:0] add_ln703_314_fu_2167_p2;
wire   [15:0] sub_ln703_170_fu_1859_p2;
wire   [15:0] add_ln703_327_fu_2204_p2;
wire   [15:0] add_ln703_325_fu_2199_p2;
wire   [15:0] add_ln703_317_fu_2182_p2;
wire   [15:0] sub_ln703_175_fu_1881_p2;
wire   [15:0] add_ln703_330_fu_2219_p2;
wire   [15:0] add_ln703_296_fu_2238_p2;
wire   [15:0] add_ln703_298_fu_2242_p2;
wire   [15:0] sub_ln703_199_fu_2246_p2;
wire   [15:0] add_ln703_301_fu_2250_p2;
wire   [15:0] add_ln703_305_fu_2254_p2;
wire   [15:0] sub_ln703_201_fu_2258_p2;
wire   [15:0] sub_ln703_205_fu_2262_p2;
wire   [15:0] sub_ln703_206_fu_2266_p2;
wire   [15:0] add_ln703_312_fu_2270_p2;
wire   [15:0] sub_ln703_207_fu_2274_p2;
wire   [15:0] sub_ln703_211_fu_2278_p2;
wire   [15:0] sub_ln703_213_fu_2282_p2;
wire   [15:0] sub_ln703_215_fu_2292_p2;
wire   [15:0] sub_ln703_216_fu_2296_p2;
wire   [15:0] add_ln703_315_fu_2300_p2;
wire   [15:0] sub_ln703_217_fu_2305_p2;
wire   [15:0] sub_ln703_218_fu_2310_p2;
wire   [15:0] sub_ln703_220_fu_2318_p2;
wire   [15:0] add_ln703_318_fu_2323_p2;
wire   [15:0] add_ln703_319_fu_2328_p2;
wire   [15:0] sub_ln703_221_fu_2332_p2;
wire   [15:0] add_ln703_320_fu_2336_p2;
wire   [15:0] sub_ln703_222_fu_2340_p2;
wire   [15:0] sub_ln703_224_fu_2348_p2;
wire   [15:0] add_ln703_321_fu_2353_p2;
wire   [15:0] sub_ln703_225_fu_2358_p2;
wire   [15:0] sub_ln703_227_fu_2368_p2;
wire   [15:0] sub_ln703_228_fu_2372_p2;
wire   [15:0] sub_ln703_229_fu_2376_p2;
wire   [15:0] sub_ln703_231_fu_2381_p2;
wire   [15:0] sub_ln703_232_fu_2385_p2;
wire   [15:0] sub_ln703_235_fu_2400_p2;
wire   [15:0] add_ln703_324_fu_2405_p2;
wire   [15:0] add_ln703_329_fu_2410_p2;
wire   [15:0] sub_ln703_219_fu_2314_p2;
wire   [15:0] sub_ln703_236_fu_2415_p2;
wire   [15:0] add_ln703_335_fu_2420_p2;
wire   [15:0] sub_ln703_238_fu_2424_p2;
wire   [15:0] sub_ln703_239_fu_2429_p2;
wire   [15:0] sub_ln703_240_fu_2434_p2;
wire   [15:0] sub_ln703_241_fu_2439_p2;
wire   [15:0] sub_ln703_242_fu_2444_p2;
wire   [15:0] sub_ln703_223_fu_2344_p2;
wire   [15:0] add_ln703_336_fu_2449_p2;
wire   [15:0] sub_ln703_243_fu_2454_p2;
wire   [15:0] add_ln703_337_fu_2459_p2;
wire   [15:0] add_ln703_339_fu_2464_p2;
wire   [15:0] sub_ln703_244_fu_2468_p2;
wire   [15:0] add_ln703_349_fu_2598_p2;
wire   [15:0] add_ln703_347_fu_2594_p2;
wire   [15:0] sub_ln703_245_fu_2472_p2;
wire   [15:0] sub_ln703_247_fu_2482_p2;
wire   [15:0] sub_ln703_248_fu_2487_p2;
wire   [15:0] add_ln703_340_fu_2491_p2;
wire   [15:0] sub_ln703_252_fu_2511_p2;
wire   [15:0] sub_ln703_253_fu_2515_p2;
wire   [15:0] sub_ln703_255_fu_2530_p2;
wire   [15:0] sub_ln703_258_fu_2544_p2;
wire   [15:0] sub_ln703_259_fu_2549_p2;
wire   [15:0] add_ln703_343_fu_2554_p2;
wire   [15:0] add_ln703_345_fu_2564_p2;
wire   [15:0] sub_ln703_226_fu_2363_p2;
wire   [15:0] add_ln703_358_fu_2672_p2;
wire   [15:0] sub_ln703_264_fu_2584_p2;
wire   [15:0] add_ln703_351_fu_2608_p2;
wire   [15:0] sub_ln703_266_fu_2618_p2;
wire   [15:0] sub_ln703_267_fu_2623_p2;
wire   [15:0] add_ln703_355_fu_2642_p2;
wire   [15:0] sub_ln703_276_fu_2667_p2;
wire   [15:0] add_ln703_361_fu_2683_p2;
wire   [15:0] sub_ln703_283_fu_2693_p2;
wire   [15:0] sub_ln703_233_fu_2390_p2;
wire   [15:0] add_ln703_370_fu_2728_p2;
wire   [15:0] add_ln703_368_fu_2723_p2;
wire   [15:0] sub_ln703_260_fu_2559_p2;
wire   [15:0] sub_ln703_214_fu_2287_p2;
wire   [15:0] add_ln703_398_fu_2747_p2;
wire   [15:0] add_ln703_523_fu_2770_p2;
wire   [15:0] sub_ln703_268_fu_2783_p2;
wire   [15:0] sub_ln703_269_fu_2787_p2;
wire   [15:0] sub_ln703_271_fu_2791_p2;
wire   [15:0] add_ln703_353_fu_2795_p2;
wire   [15:0] add_ln703_357_fu_2811_p2;
wire   [15:0] sub_ln703_279_fu_2815_p2;
wire   [15:0] sub_ln703_280_fu_2819_p2;
wire   [15:0] add_ln703_363_fu_2823_p2;
wire   [15:0] add_ln703_364_fu_2831_p2;
wire   [15:0] sub_ln703_285_fu_2836_p2;
wire   [15:0] add_ln703_365_fu_2841_p2;
wire   [15:0] sub_ln703_286_fu_2845_p2;
wire   [15:0] sub_ln703_290_fu_2859_p2;
wire   [15:0] sub_ln703_273_fu_2799_p2;
wire   [15:0] sub_ln703_291_fu_2863_p2;
wire   [15:0] sub_ln703_292_fu_2867_p2;
wire   [15:0] add_ln703_366_fu_2871_p2;
wire   [15:0] sub_ln703_295_fu_2880_p2;
wire   [15:0] sub_ln703_297_fu_2884_p2;
wire   [15:0] sub_ln703_298_fu_2889_p2;
wire   [15:0] sub_ln703_299_fu_2894_p2;
wire   [15:0] sub_ln703_300_fu_2898_p2;
wire   [15:0] add_ln703_367_fu_2903_p2;
wire   [15:0] sub_ln703_302_fu_2907_p2;
wire   [15:0] add_ln703_385_fu_3011_p2;
wire   [15:0] add_ln703_383_fu_3007_p2;
wire   [15:0] sub_ln703_303_fu_2912_p2;
wire   [15:0] sub_ln703_304_fu_2917_p2;
wire   [15:0] add_ln703_372_fu_2927_p2;
wire   [15:0] sub_ln703_306_fu_2931_p2;
wire   [15:0] add_ln703_374_fu_2936_p2;
wire   [15:0] add_ln703_387_fu_3046_p2;
wire   [15:0] sub_ln703_307_fu_2941_p2;
wire   [15:0] sub_ln703_308_fu_2946_p2;
wire   [15:0] sub_ln703_309_fu_2951_p2;
wire   [15:0] add_ln703_377_fu_2956_p2;
wire   [15:0] add_ln703_378_fu_2960_p2;
wire   [15:0] sub_ln703_277_fu_2803_p2;
wire   [15:0] add_ln703_392_fu_3081_p2;
wire   [15:0] add_ln703_379_fu_2964_p2;
wire   [15:0] add_ln703_380_fu_2969_p2;
wire   [15:0] add_ln703_381_fu_2973_p2;
wire   [15:0] add_ln703_382_fu_2983_p2;
wire   [15:0] sub_ln703_311_fu_2988_p2;
wire   [15:0] sub_ln703_282_fu_2827_p2;
wire   [15:0] add_ln703_395_fu_3116_p2;
wire   [15:0] sub_ln703_312_fu_2993_p2;
wire   [15:0] add_ln703_403_fu_3131_p2;
wire   [15:0] sub_ln703_314_fu_3003_p2;
wire   [15:0] add_ln703_406_fu_3145_p2;
wire   [15:0] sub_ln703_316_fu_3026_p2;
wire   [15:0] sub_ln703_305_fu_2922_p2;
wire   [15:0] sub_ln703_288_fu_2854_p2;
wire   [15:0] add_ln703_414_fu_3165_p2;
wire   [15:0] sub_ln703_318_fu_3036_p2;
wire   [15:0] add_ln703_391_fu_3061_p2;
wire   [15:0] sub_ln703_321_fu_3066_p2;
wire   [15:0] sub_ln703_322_fu_3071_p2;
wire   [15:0] sub_ln703_323_fu_3076_p2;
wire   [15:0] add_ln703_394_fu_3086_p2;
wire   [15:0] sub_ln703_324_fu_3091_p2;
wire   [15:0] sub_ln703_325_fu_3096_p2;
wire   [15:0] sub_ln703_327_fu_3106_p2;
wire   [15:0] add_ln703_397_fu_3121_p2;
wire   [15:0] add_ln703_419_fu_3225_p2;
wire   [15:0] add_ln703_404_fu_3135_p2;
wire   [15:0] sub_ln703_331_fu_3140_p2;
wire   [15:0] add_ln703_413_fu_3160_p2;
wire   [15:0] sub_ln703_287_fu_2849_p2;
wire   [15:0] add_ln703_425_fu_3254_p2;
wire   [15:0] add_ln703_423_fu_3249_p2;
wire   [15:0] sub_ln703_317_fu_3031_p2;
wire   [15:0] sub_ln703_337_fu_3190_p2;
wire   [15:0] sub_ln703_338_fu_3195_p2;
wire   [15:0] sub_ln703_294_fu_2875_p2;
wire   [15:0] add_ln703_432_fu_3279_p2;
wire   [15:0] add_ln703_418_fu_3210_p2;
wire   [15:0] add_ln703_421_fu_3229_p2;
wire   [15:0] add_ln703_422_fu_3239_p2;
wire   [15:0] add_ln703_428_fu_3264_p2;
wire   [15:0] sub_ln703_320_fu_3056_p2;
wire   [15:0] sub_ln703_310_fu_2978_p2;
wire   [15:0] sub_ln703_357_fu_3295_p2;
wire   [15:0] sub_ln703_319_fu_3041_p2;
wire   [15:0] sub_ln703_329_fu_3126_p2;
wire   [15:0] sub_ln703_278_fu_2807_p2;
wire   [15:0] sub_ln703_332_fu_3376_p2;
wire   [15:0] add_ln703_411_fu_3380_p2;
wire   [15:0] sub_ln703_335_fu_3384_p2;
wire   [15:0] sub_ln703_346_fu_3396_p2;
wire   [15:0] sub_ln703_349_fu_3410_p2;
wire   [15:0] add_ln703_429_fu_3418_p2;
wire   [15:0] add_ln703_430_fu_3423_p2;
wire   [15:0] sub_ln703_352_fu_3427_p2;
wire   [15:0] sub_ln703_354_fu_3431_p2;
wire   [15:0] sub_ln703_355_fu_3435_p2;
wire   [15:0] sub_ln703_341_fu_3388_p2;
wire   [15:0] add_ln703_436_fu_3439_p2;
wire   [15:0] add_ln703_437_fu_3443_p2;
wire   [15:0] sub_ln703_348_fu_3405_p2;
wire   [15:0] sub_ln703_359_fu_3448_p2;
wire   [15:0] sub_ln703_360_fu_3453_p2;
wire   [15:0] sub_ln703_351_fu_3414_p2;
wire   [15:0] add_ln703_459_fu_3557_p2;
wire   [15:0] add_ln703_440_fu_3466_p2;
wire   [15:0] sub_ln703_364_fu_3470_p2;
wire   [15:0] add_ln703_441_fu_3480_p2;
wire   [15:0] sub_ln703_366_fu_3484_p2;
wire   [15:0] sub_ln703_367_fu_3488_p2;
wire   [15:0] sub_ln703_368_fu_3493_p2;
wire   [15:0] sub_ln703_369_fu_3497_p2;
wire   [15:0] add_ln703_442_fu_3502_p2;
wire   [15:0] add_ln703_444_fu_3506_p2;
wire   [15:0] add_ln703_448_fu_3511_p2;
wire   [15:0] sub_ln703_370_fu_3515_p2;
wire   [15:0] add_ln703_450_fu_3520_p2;
wire   [15:0] sub_ln703_330_fu_3372_p2;
wire   [15:0] add_ln703_467_fu_3635_p2;
wire   [15:0] add_ln703_465_fu_3630_p2;
wire   [15:0] add_ln703_452_fu_3524_p2;
wire   [15:0] add_ln703_453_fu_3528_p2;
wire   [15:0] sub_ln703_372_fu_3532_p2;
wire   [15:0] add_ln703_455_fu_3537_p2;
wire   [15:0] add_ln703_456_fu_3542_p2;
wire   [15:0] add_ln703_458_fu_3552_p2;
wire   [15:0] add_ln703_461_fu_3561_p2;
wire   [15:0] sub_ln703_363_fu_3461_p2;
wire   [15:0] add_ln703_462_fu_3571_p2;
wire   [15:0] sub_ln703_375_fu_3576_p2;
wire   [15:0] add_ln703_463_fu_3581_p2;
wire   [15:0] add_ln703_464_fu_3586_p2;
wire   [15:0] sub_ln703_377_fu_3596_p2;
wire   [15:0] sub_ln703_378_fu_3601_p2;
wire   [15:0] sub_ln703_379_fu_3606_p2;
wire   [15:0] sub_ln703_380_fu_3611_p2;
wire   [15:0] sub_ln703_381_fu_3616_p2;
wire   [15:0] sub_ln703_343_fu_3392_p2;
wire   [15:0] add_ln703_479_fu_3735_p2;
wire   [15:0] sub_ln703_382_fu_3621_p2;
wire   [15:0] sub_ln703_383_fu_3626_p2;
wire   [15:0] add_ln703_468_fu_3639_p2;
wire   [15:0] sub_ln703_385_fu_3650_p2;
wire   [15:0] sub_ln703_361_fu_3457_p2;
wire   [15:0] add_ln703_489_fu_3771_p2;
wire   [15:0] sub_ln703_388_fu_3670_p2;
wire   [15:0] sub_ln703_389_fu_3675_p2;
wire   [15:0] add_ln703_474_fu_3680_p2;
wire   [15:0] sub_ln703_374_fu_3566_p2;
wire   [15:0] sub_ln703_365_fu_3475_p2;
wire   [15:0] add_ln703_494_fu_3801_p2;
wire   [15:0] sub_ln703_391_fu_3695_p2;
wire   [15:0] sub_ln703_392_fu_3700_p2;
wire   [15:0] add_ln703_500_fu_3821_p2;
wire   [15:0] add_ln703_504_fu_3830_p2;
wire   [15:0] add_ln703_505_fu_3834_p2;
wire   [15:0] add_ln703_501_fu_3825_p2;
wire   [15:0] add_ln703_477_fu_3715_p2;
wire   [15:0] add_ln703_482_fu_3740_p2;
wire   [15:0] add_ln703_487_fu_3756_p2;
wire   [15:0] add_ln703_488_fu_3766_p2;
wire   [15:0] add_ln703_491_fu_3776_p2;
wire   [15:0] add_ln703_511_fu_3874_p2;
wire   [15:0] add_ln703_509_fu_3870_p2;
wire   [15:0] add_ln703_493_fu_3796_p2;
wire   [15:0] sub_ln703_396_fu_3725_p2;
wire   [15:0] sub_ln703_397_fu_3746_p2;
wire   [15:0] sub_ln703_398_fu_3751_p2;
wire   [15:0] add_ln703_536_fu_3908_p2;
wire   [15:0] add_ln703_532_fu_3904_p2;
wire   [15:0] sub_ln703_373_fu_3547_p2;
wire   [15:0] add_ln703_542_fu_3918_p2;
wire   [15:0] sub_ln703_376_fu_3591_p2;
wire   [15:0] add_ln703_553_fu_3928_p2;
wire   [15:0] add_ln703_519_fu_3899_p2;
wire   [15:0] sub_ln703_347_fu_3400_p2;
wire   [15:0] add_ln703_564_fu_3947_p2;
wire   [15:0] sub_ln703_400_fu_3973_p2;
wire   [15:0] sub_ln703_404_fu_3977_p2;
wire   [15:0] sub_ln703_407_fu_3985_p2;
wire   [15:0] sub_ln703_409_fu_3989_p2;
wire   [15:0] sub_ln703_410_fu_3993_p2;
wire   [15:0] sub_ln703_413_fu_3997_p2;
wire   [15:0] add_ln703_529_fu_4071_p2;
wire   [15:0] add_ln703_508_fu_4006_p2;
wire   [15:0] add_ln703_539_fu_4085_p2;
wire   [15:0] sub_ln703_417_fu_4010_p2;
wire   [15:0] sub_ln703_418_fu_4014_p2;
wire   [15:0] sub_ln703_420_fu_4019_p2;
wire   [15:0] sub_ln703_421_fu_4023_p2;
wire   [15:0] sub_ln703_422_fu_4027_p2;
wire   [15:0] sub_ln703_423_fu_4031_p2;
wire   [15:0] add_ln703_513_fu_4035_p2;
wire   [15:0] sub_ln703_424_fu_4040_p2;
wire   [15:0] sub_ln703_426_fu_4049_p2;
wire   [15:0] sub_ln703_427_fu_4054_p2;
wire   [15:0] add_ln703_520_fu_4058_p2;
wire   [15:0] add_ln703_521_fu_4062_p2;
wire   [15:0] add_ln703_522_fu_4067_p2;
wire   [15:0] add_ln703_538_fu_4075_p2;
wire   [15:0] sub_ln703_428_fu_4080_p2;
wire   [15:0] add_ln703_541_fu_4089_p2;
wire   [15:0] add_ln703_546_fu_4094_p2;
wire   [15:0] add_ln703_548_fu_4098_p2;
wire   [15:0] sub_ln703_429_fu_4102_p2;
wire   [15:0] sub_ln703_430_fu_4106_p2;
wire   [15:0] add_ln703_550_fu_4111_p2;
wire   [15:0] add_ln703_551_fu_4115_p2;
wire   [15:0] sub_ln703_431_fu_4120_p2;
wire   [15:0] sub_ln703_432_fu_4124_p2;
wire   [15:0] add_ln703_552_fu_4139_p2;
wire   [15:0] sub_ln703_436_fu_4149_p2;
wire   [15:0] sub_ln703_425_fu_4044_p2;
wire   [15:0] sub_ln703_437_fu_4154_p2;
wire   [15:0] add_ln703_557_fu_4158_p2;
wire   [15:0] sub_ln703_439_fu_4168_p2;
wire   [15:0] sub_ln703_441_fu_4172_p2;
wire   [15:0] sub_ln703_443_fu_4182_p2;
wire   [15:0] add_ln703_570_fu_4294_p2;
wire   [15:0] sub_ln703_445_fu_4192_p2;
wire   [15:0] sub_ln703_446_fu_4197_p2;
wire   [15:0] sub_ln703_447_fu_4202_p2;
wire   [15:0] add_ln703_558_fu_4216_p2;
wire   [15:0] sub_ln703_450_fu_4221_p2;
wire   [15:0] sub_ln703_451_fu_4226_p2;
wire   [15:0] add_ln703_559_fu_4241_p2;
wire   [15:0] sub_ln703_433_fu_4129_p2;
wire   [15:0] sub_ln703_406_fu_3981_p2;
wire   [15:0] add_ln703_577_fu_4343_p2;
wire   [15:0] sub_ln703_454_fu_4246_p2;
wire   [15:0] sub_ln703_455_fu_4251_p2;
wire   [15:0] sub_ln703_435_fu_4144_p2;
wire   [15:0] sub_ln703_456_fu_4255_p2;
wire   [15:0] add_ln703_561_fu_4260_p2;
wire   [15:0] sub_ln703_457_fu_4265_p2;
wire   [15:0] sub_ln703_438_fu_4163_p2;
wire   [15:0] add_ln703_562_fu_4275_p2;
wire   [15:0] add_ln703_563_fu_4280_p2;
wire   [15:0] sub_ln703_460_fu_4289_p2;
wire   [15:0] sub_ln703_415_fu_4001_p2;
wire   [15:0] add_ln703_589_fu_4408_p2;
wire   [15:0] add_ln703_587_fu_4403_p2;
wire   [15:0] add_ln703_571_fu_4298_p2;
wire   [15:0] sub_ln703_464_fu_4318_p2;
wire   [15:0] sub_ln703_465_fu_4328_p2;
wire   [15:0] add_ln703_597_fu_4437_p2;
wire   [15:0] add_ln703_594_fu_4433_p2;
wire   [15:0] add_ln703_576_fu_4338_p2;
wire   [15:0] add_ln703_580_fu_4348_p2;
wire   [15:0] sub_ln703_471_fu_4378_p2;
wire   [15:0] add_ln703_585_fu_4383_p2;
wire   [15:0] sub_ln703_473_fu_4388_p2;
wire   [15:0] sub_ln703_474_fu_4393_p2;
wire   [15:0] sub_ln703_442_fu_4177_p2;
wire   [15:0] add_ln703_602_fu_4482_p2;
wire   [15:0] add_ln703_607_fu_4491_p2;
wire   [15:0] add_ln703_604_fu_4486_p2;
wire   [15:0] sub_ln703_444_fu_4187_p2;
wire   [15:0] sub_ln703_449_fu_4211_p2;
wire   [15:0] add_ln703_614_fu_4506_p2;
wire   [15:0] sub_ln703_492_fu_4472_p2;
wire   [15:0] add_ln703_608_fu_4495_p2;
wire   [15:0] sub_ln703_434_fu_4134_p2;
wire   [15:0] add_ln703_631_fu_4526_p2;
wire   [15:0] sub_ln703_459_fu_4284_p2;
wire   [15:0] add_ln703_574_fu_4566_p2;
wire   [15:0] sub_ln703_472_fu_4570_p2;
wire   [15:0] sub_ln703_477_fu_4578_p2;
wire   [15:0] sub_ln703_478_fu_4582_p2;
wire   [15:0] sub_ln703_479_fu_4586_p2;
wire   [15:0] sub_ln703_480_fu_4590_p2;
wire   [15:0] sub_ln703_481_fu_4595_p2;
wire   [15:0] sub_ln703_484_fu_4599_p2;
wire   [15:0] sub_ln703_485_fu_4603_p2;
wire   [15:0] sub_ln703_486_fu_4607_p2;
wire   [15:0] add_ln703_601_fu_4620_p2;
wire   [15:0] sub_ln703_493_fu_4624_p2;
wire   [15:0] add_ln703_611_fu_4628_p2;
wire   [15:0] sub_ln703_494_fu_4632_p2;
wire   [15:0] sub_ln703_476_fu_4574_p2;
wire   [15:0] add_ln703_612_fu_4640_p2;
wire   [15:0] add_ln703_613_fu_4645_p2;
wire   [15:0] sub_ln703_496_fu_4650_p2;
wire   [15:0] sub_ln703_497_fu_4654_p2;
wire   [15:0] sub_ln703_498_fu_4659_p2;
wire   [15:0] sub_ln703_466_fu_4562_p2;
wire   [15:0] add_ln703_624_fu_4754_p2;
wire   [15:0] sub_ln703_500_fu_4668_p2;
wire   [15:0] sub_ln703_501_fu_4672_p2;
wire   [15:0] add_ln703_617_fu_4677_p2;
wire   [15:0] sub_ln703_502_fu_4682_p2;
wire   [15:0] add_ln703_618_fu_4687_p2;
wire   [15:0] sub_ln703_487_fu_4611_p2;
wire   [15:0] add_ln703_619_fu_4692_p2;
wire   [15:0] sub_ln703_489_fu_4615_p2;
wire   [15:0] add_ln703_620_fu_4696_p2;
wire   [15:0] sub_ln703_504_fu_4700_p2;
wire   [15:0] sub_ln703_506_fu_4705_p2;
wire   [15:0] sub_ln703_507_fu_4710_p2;
wire   [15:0] sub_ln703_508_fu_4715_p2;
wire   [15:0] add_ln703_622_fu_4720_p2;
wire   [15:0] sub_ln703_511_fu_4735_p2;
wire   [15:0] add_ln703_623_fu_4739_p2;
wire   [15:0] sub_ln703_512_fu_4744_p2;
wire   [15:0] add_ln703_626_fu_4759_p2;
wire   [15:0] sub_ln703_499_fu_4663_p2;
wire   [15:0] sub_ln703_514_fu_4764_p2;
wire   [15:0] add_ln703_627_fu_4769_p2;
wire   [15:0] add_ln703_629_fu_4774_p2;
wire   [15:0] sub_ln703_515_fu_4778_p2;
wire   [15:0] sub_ln703_516_fu_4783_p2;
wire   [15:0] sub_ln703_517_fu_4788_p2;
wire   [15:0] add_ln703_636_fu_4793_p2;
wire   [15:0] sub_ln703_518_fu_4798_p2;
wire   [15:0] add_ln703_638_fu_4803_p2;
wire   [15:0] sub_ln703_520_fu_4813_p2;
wire   [15:0] add_ln703_642_fu_4817_p2;
wire   [15:0] add_ln703_643_fu_4821_p2;
wire   [15:0] add_ln703_644_fu_4826_p2;
wire   [15:0] add_ln703_645_fu_4835_p2;
wire   [15:0] sub_ln703_522_fu_4840_p2;
wire   [15:0] sub_ln703_523_fu_4845_p2;
wire   [15:0] sub_ln703_510_fu_4730_p2;
wire   [15:0] sub_ln703_463_fu_4558_p2;
wire   [15:0] add_ln703_655_fu_4969_p2;
wire   [15:0] add_ln703_653_fu_4964_p2;
wire   [15:0] sub_ln703_524_fu_4850_p2;
wire   [15:0] sub_ln703_525_fu_4855_p2;
wire   [15:0] sub_ln703_513_fu_4749_p2;
wire   [15:0] sub_ln703_531_fu_4890_p2;
wire   [15:0] sub_ln703_534_fu_4909_p2;
wire   [15:0] add_ln703_649_fu_4914_p2;
wire   [15:0] add_ln703_663_fu_5009_p2;
wire   [15:0] sub_ln703_521_fu_4830_p2;
wire   [15:0] add_ln703_656_fu_4973_p2;
wire   [15:0] sub_ln703_543_fu_4979_p2;
wire   [15:0] add_ln703_658_fu_4989_p2;
wire   [15:0] sub_ln703_530_fu_4885_p2;
wire   [15:0] add_ln703_675_fu_5048_p2;
wire   [15:0] add_ln703_673_fu_5044_p2;
wire   [15:0] add_ln703_681_fu_5062_p2;
wire   [15:0] add_ln703_678_fu_5058_p2;
wire   [15:0] sub_ln703_519_fu_4808_p2;
wire   [15:0] add_ln703_683_fu_5072_p2;
wire   [15:0] sub_ln703_536_fu_4924_p2;
wire   [15:0] sub_ln703_537_fu_4929_p2;
wire   [15:0] sub_ln703_528_fu_4875_p2;
wire   [15:0] add_ln703_671_fu_5039_p2;
wire   [15:0] add_ln703_687_fu_5082_p2;
wire   [15:0] add_ln703_689_fu_5087_p2;
wire   [15:0] sub_ln703_509_fu_4725_p2;
wire   [15:0] sub_ln703_495_fu_4636_p2;
wire   [15:0] sub_ln703_546_fu_5142_p2;
wire   [15:0] sub_ln703_547_fu_5146_p2;
wire   [15:0] add_ln703_659_fu_5150_p2;
wire   [15:0] sub_ln703_548_fu_5154_p2;
wire   [15:0] sub_ln703_550_fu_5162_p2;
wire   [15:0] add_ln703_662_fu_5166_p2;
wire   [15:0] sub_ln703_553_fu_5174_p2;
wire   [15:0] sub_ln703_554_fu_5178_p2;
wire   [15:0] sub_ln703_555_fu_5182_p2;
wire   [15:0] add_ln703_669_fu_5186_p2;
wire   [15:0] sub_ln703_560_fu_5195_p2;
wire   [15:0] sub_ln703_561_fu_5200_p2;
wire   [15:0] sub_ln703_562_fu_5205_p2;
wire   [15:0] sub_ln703_564_fu_5214_p2;
wire   [15:0] sub_ln703_565_fu_5219_p2;
wire   [15:0] sub_ln703_566_fu_5223_p2;
wire   [15:0] sub_ln703_567_fu_5227_p2;
wire   [15:0] sub_ln703_568_fu_5232_p2;
wire   [15:0] add_ln703_702_fu_5332_p2;
wire   [15:0] sub_ln703_569_fu_5236_p2;
wire   [15:0] add_ln703_690_fu_5240_p2;
wire   [15:0] add_ln703_692_fu_5245_p2;
wire   [15:0] add_ln703_693_fu_5249_p2;
wire   [15:0] add_ln703_708_fu_5361_p2;
wire   [15:0] add_ln703_694_fu_5254_p2;
wire   [15:0] add_ln703_695_fu_5259_p2;
wire   [15:0] sub_ln703_570_fu_5263_p2;
wire   [15:0] sub_ln703_571_fu_5267_p2;
wire   [15:0] sub_ln703_545_fu_5138_p2;
wire   [15:0] add_ln703_710_fu_5390_p2;
wire   [15:0] add_ln703_696_fu_5272_p2;
wire   [15:0] sub_ln703_559_fu_5190_p2;
wire   [15:0] sub_ln703_572_fu_5276_p2;
wire   [15:0] add_ln703_699_fu_5281_p2;
wire   [15:0] add_ln703_700_fu_5285_p2;
wire   [15:0] sub_ln703_574_fu_5290_p2;
wire   [15:0] sub_ln703_563_fu_5209_p2;
wire   [15:0] sub_ln703_576_fu_5299_p2;
wire   [15:0] sub_ln703_577_fu_5304_p2;
wire   [15:0] add_ln703_701_fu_5313_p2;
wire   [15:0] sub_ln703_579_fu_5318_p2;
wire   [15:0] sub_ln703_580_fu_5323_p2;
wire   [15:0] sub_ln703_581_fu_5328_p2;
wire   [15:0] add_ln703_727_fu_5481_p2;
wire   [15:0] add_ln703_724_fu_5477_p2;
wire   [15:0] sub_ln703_587_fu_5356_p2;
wire   [15:0] add_ln703_709_fu_5365_p2;
wire   [15:0] sub_ln703_588_fu_5370_p2;
wire   [15:0] sub_ln703_590_fu_5380_p2;
wire   [15:0] sub_ln703_591_fu_5385_p2;
wire   [15:0] add_ln703_712_fu_5395_p2;
wire   [15:0] add_ln703_714_fu_5405_p2;
wire   [15:0] add_ln703_715_fu_5425_p2;
wire   [15:0] add_ln703_716_fu_5429_p2;
wire   [15:0] add_ln703_718_fu_5434_p2;
wire   [15:0] sub_ln703_596_fu_5444_p2;
wire   [15:0] sub_ln703_578_fu_5308_p2;
wire   [15:0] sub_ln703_597_fu_5449_p2;
wire   [15:0] sub_ln703_599_fu_5459_p2;
wire   [15:0] sub_ln703_600_fu_5464_p2;
wire   [15:0] add_ln703_720_fu_5469_p2;
wire   [15:0] sub_ln703_601_fu_5473_p2;
wire   [15:0] sub_ln703_552_fu_5170_p2;
wire   [15:0] add_ln703_738_fu_5581_p2;
wire   [15:0] add_ln703_736_fu_5576_p2;
wire   [15:0] sub_ln703_584_fu_5341_p2;
wire   [15:0] sub_ln703_607_fu_5506_p2;
wire   [15:0] sub_ln703_592_fu_5400_p2;
wire   [15:0] sub_ln703_575_fu_5295_p2;
wire   [15:0] add_ln703_745_fu_5606_p2;
wire   [15:0] sub_ln703_549_fu_5158_p2;
wire   [15:0] add_ln703_750_fu_5616_p2;
wire   [15:0] add_ln703_730_fu_5541_p2;
wire   [15:0] add_ln703_732_fu_5546_p2;
wire   [15:0] sub_ln703_617_fu_5561_p2;
wire   [15:0] add_ln703_739_fu_5585_p2;
wire   [15:0] add_ln703_741_fu_5591_p2;
wire   [15:0] add_ln703_744_fu_5601_p2;
wire   [15:0] add_ln703_747_fu_5611_p2;
wire   [15:0] add_ln703_753_fu_5621_p2;
wire   [15:0] sub_ln703_585_fu_5346_p2;
wire   [15:0] sub_ln703_602_fu_5688_p2;
wire   [15:0] add_ln703_721_fu_5692_p2;
wire   [15:0] add_ln703_729_fu_5700_p2;
wire   [15:0] sub_ln703_615_fu_5708_p2;
wire   [15:0] sub_ln703_619_fu_5716_p2;
wire   [15:0] sub_ln703_620_fu_5721_p2;
wire   [15:0] sub_ln703_622_fu_5730_p2;
wire   [15:0] sub_ln703_623_fu_5734_p2;
wire   [15:0] add_ln703_742_fu_5738_p2;
wire   [15:0] sub_ln703_606_fu_5696_p2;
wire   [15:0] sub_ln703_625_fu_5742_p2;
wire   [15:0] sub_ln703_626_fu_5746_p2;
wire   [15:0] sub_ln703_627_fu_5750_p2;
wire   [15:0] sub_ln703_611_fu_5704_p2;
wire   [15:0] sub_ln703_628_fu_5755_p2;
wire   [15:0] add_ln703_748_fu_5759_p2;
wire   [15:0] sub_ln703_629_fu_5763_p2;
wire   [15:0] sub_ln703_632_fu_5768_p2;
wire   [15:0] sub_ln703_633_fu_5772_p2;
wire   [15:0] add_ln703_754_fu_5776_p2;
wire   [15:0] sub_ln703_635_fu_5780_p2;
wire   [15:0] sub_ln703_621_fu_5726_p2;
wire   [15:0] sub_ln703_640_fu_5794_p2;
wire   [15:0] sub_ln703_642_fu_5804_p2;
wire   [15:0] add_ln703_756_fu_5809_p2;
wire   [15:0] add_ln703_757_fu_5814_p2;
wire   [15:0] add_ln703_759_fu_5818_p2;
wire   [15:0] sub_ln703_643_fu_5822_p2;
wire   [15:0] sub_ln703_646_fu_5832_p2;
wire   [15:0] add_ln703_761_fu_5837_p2;
wire   [15:0] add_ln703_769_fu_5946_p2;
wire   [15:0] add_ln703_767_fu_5942_p2;
wire   [15:0] add_ln703_763_fu_5842_p2;
wire   [15:0] sub_ln703_647_fu_5846_p2;
wire   [15:0] sub_ln703_649_fu_5851_p2;
wire   [15:0] sub_ln703_651_fu_5856_p2;
wire   [15:0] add_ln703_764_fu_5861_p2;
wire   [15:0] sub_ln703_652_fu_5865_p2;
wire   [15:0] sub_ln703_616_fu_5712_p2;
wire   [15:0] add_ln703_775_fu_5994_p2;
wire   [15:0] sub_ln703_653_fu_5870_p2;
wire   [15:0] sub_ln703_654_fu_5875_p2;
wire   [15:0] sub_ln703_655_fu_5879_p2;
wire   [15:0] sub_ln703_656_fu_5884_p2;
wire   [15:0] sub_ln703_636_fu_5784_p2;
wire   [15:0] sub_ln703_657_fu_5889_p2;
wire   [15:0] add_ln703_785_fu_6038_p2;
wire   [15:0] add_ln703_766_fu_5893_p2;
wire   [15:0] sub_ln703_658_fu_5898_p2;
wire   [15:0] sub_ln703_659_fu_5903_p2;
wire   [15:0] sub_ln703_660_fu_5908_p2;
wire   [15:0] sub_ln703_664_fu_5928_p2;
wire   [15:0] sub_ln703_666_fu_5937_p2;
wire   [15:0] add_ln703_771_fu_5961_p2;
wire   [15:0] add_ln703_772_fu_5966_p2;
wire   [15:0] sub_ln703_668_fu_5971_p2;
wire   [15:0] sub_ln703_670_fu_5980_p2;
wire   [15:0] add_ln703_774_fu_5985_p2;
wire   [15:0] sub_ln703_671_fu_5989_p2;
wire   [15:0] add_ln703_777_fu_5999_p2;
wire   [15:0] sub_ln703_672_fu_6004_p2;
wire   [15:0] sub_ln703_673_fu_6009_p2;
wire   [15:0] sub_ln703_674_fu_6014_p2;
wire   [15:0] sub_ln703_675_fu_6019_p2;
wire   [15:0] add_ln703_781_fu_6029_p2;
wire   [15:0] add_ln703_786_fu_6042_p2;
wire   [15:0] sub_ln703_677_fu_6047_p2;
wire   [15:0] sub_ln703_641_fu_5799_p2;
wire   [15:0] add_ln703_795_fu_6156_p2;
wire   [15:0] add_ln703_794_fu_6151_p2;
wire   [15:0] sub_ln703_663_fu_5923_p2;
wire   [15:0] add_ln703_788_fu_6082_p2;
wire   [15:0] sub_ln703_689_fu_6096_p2;
wire   [15:0] add_ln703_790_fu_6121_p2;
wire   [15:0] sub_ln703_639_fu_5789_p2;
wire   [15:0] sub_ln703_661_fu_5913_p2;
wire   [15:0] add_ln703_817_fu_6201_p2;
wire   [15:0] add_ln703_815_fu_6196_p2;
wire   [15:0] sub_ln703_645_fu_5827_p2;
wire   [15:0] add_ln703_820_fu_6211_p2;
wire   [15:0] sub_ln703_681_fu_6238_p2;
wire   [15:0] sub_ln703_683_fu_6242_p2;
wire   [15:0] sub_ln703_685_fu_6246_p2;
wire   [15:0] add_ln703_789_fu_6250_p2;
wire   [15:0] sub_ln703_695_fu_6254_p2;
wire   [15:0] add_ln703_803_fu_6319_p2;
wire   [15:0] add_ln703_793_fu_6258_p2;
wire   [15:0] add_ln703_797_fu_6262_p2;
wire   [15:0] sub_ln703_698_fu_6267_p2;
wire   [15:0] sub_ln703_699_fu_6271_p2;
wire   [15:0] add_ln703_799_fu_6276_p2;
wire   [15:0] add_ln703_807_fu_6369_p2;
wire   [15:0] sub_ln703_701_fu_6281_p2;
wire   [15:0] sub_ln703_702_fu_6285_p2;
wire   [15:0] sub_ln703_703_fu_6289_p2;
wire   [15:0] sub_ln703_708_fu_6302_p2;
wire   [15:0] sub_ln703_709_fu_6306_p2;
wire   [15:0] add_ln703_800_fu_6315_p2;
wire   [15:0] add_ln703_804_fu_6323_p2;
wire   [15:0] sub_ln703_713_fu_6337_p2;
wire   [15:0] add_ln703_805_fu_6341_p2;
wire   [15:0] sub_ln703_714_fu_6345_p2;
wire   [15:0] sub_ln703_715_fu_6350_p2;
wire   [15:0] add_ln703_806_fu_6359_p2;
wire   [15:0] add_ln703_808_fu_6373_p2;
wire   [15:0] add_ln703_809_fu_6378_p2;
wire   [15:0] sub_ln703_718_fu_6382_p2;
wire   [15:0] sub_ln703_719_fu_6386_p2;
wire   [15:0] sub_ln703_720_fu_6391_p2;
wire   [15:0] add_ln703_810_fu_6396_p2;
wire   [15:0] add_ln703_811_fu_6401_p2;
wire   [15:0] add_ln703_812_fu_6405_p2;
wire   [15:0] add_ln703_813_fu_6409_p2;
wire   [15:0] sub_ln703_721_fu_6413_p2;
wire   [15:0] add_ln703_823_fu_6512_p2;
wire   [15:0] add_ln703_814_fu_6417_p2;
wire   [15:0] sub_ln703_722_fu_6422_p2;
wire   [15:0] sub_ln703_710_fu_6311_p2;
wire   [15:0] sub_ln703_712_fu_6332_p2;
wire   [15:0] sub_ln703_725_fu_6437_p2;
wire   [15:0] add_ln703_830_fu_6550_p2;
wire   [15:0] add_ln703_829_fu_6546_p2;
wire   [15:0] sub_ln703_726_fu_6442_p2;
wire   [15:0] add_ln703_832_fu_6569_p2;
wire   [15:0] sub_ln703_729_fu_6462_p2;
wire   [15:0] sub_ln703_730_fu_6467_p2;
wire   [15:0] sub_ln703_731_fu_6472_p2;
wire   [15:0] sub_ln703_732_fu_6477_p2;
wire   [15:0] add_ln703_822_fu_6482_p2;
wire   [15:0] sub_ln703_734_fu_6492_p2;
wire   [15:0] sub_ln703_735_fu_6497_p2;
wire   [15:0] sub_ln703_737_fu_6507_p2;
wire   [15:0] add_ln703_824_fu_6516_p2;
wire   [15:0] sub_ln703_723_fu_6427_p2;
wire   [15:0] add_ln703_828_fu_6536_p2;
wire   [15:0] sub_ln703_739_fu_6541_p2;
wire   [15:0] sub_ln703_740_fu_6560_p2;
wire   [15:0] sub_ln703_744_fu_6565_p2;
wire   [15:0] sub_ln703_747_fu_6584_p2;
wire   [15:0] sub_ln703_748_fu_6589_p2;
wire   [15:0] sub_ln703_751_fu_6604_p2;
wire   [15:0] sub_ln703_752_fu_6609_p2;
wire   [15:0] sub_ln703_705_fu_6294_p2;
wire   [15:0] add_ln703_843_fu_6674_p2;
wire   [15:0] add_ln703_842_fu_6669_p2;
wire   [15:0] sub_ln703_753_fu_6614_p2;
wire   [15:0] sub_ln703_754_fu_6619_p2;
wire   [15:0] add_ln703_850_fu_6698_p2;
wire   [15:0] add_ln703_848_fu_6694_p2;
wire   [15:0] add_ln703_837_fu_6624_p2;
wire   [15:0] sub_ln703_711_fu_6328_p2;
wire   [15:0] add_ln703_853_fu_6718_p2;
wire   [15:0] add_ln703_852_fu_6713_p2;
wire   [15:0] sub_ln703_716_fu_6354_p2;
wire   [15:0] add_ln703_857_fu_6728_p2;
wire   [15:0] add_ln703_844_fu_6678_p2;
wire   [15:0] sub_ln703_706_fu_6298_p2;
wire   [15:0] add_ln703_863_fu_6744_p2;
wire   [15:0] add_ln703_854_fu_6722_p2;
wire   [15:0] add_ln703_864_fu_6749_p2;
wire   [15:0] sub_ln703_717_fu_6364_p2;
wire   [15:0] sub_ln703_738_fu_6521_p2;
wire   [15:0] sub_ln703_741_fu_6795_p2;
wire   [15:0] sub_ln703_743_fu_6803_p2;
wire   [15:0] sub_ln703_750_fu_6811_p2;
wire   [15:0] add_ln703_835_fu_6815_p2;
wire   [15:0] sub_ln703_755_fu_6819_p2;
wire   [15:0] sub_ln703_756_fu_6823_p2;
wire   [15:0] sub_ln703_758_fu_6827_p2;
wire   [15:0] sub_ln703_760_fu_6831_p2;
wire   [15:0] sub_ln703_742_fu_6799_p2;
wire   [15:0] add_ln703_839_fu_6836_p2;
wire   [15:0] sub_ln703_745_fu_6807_p2;
wire   [15:0] sub_ln703_762_fu_6841_p2;
wire   [15:0] sub_ln703_764_fu_6845_p2;
wire   [15:0] sub_ln703_765_fu_6849_p2;
wire   [15:0] sub_ln703_766_fu_6853_p2;
wire   [15:0] add_ln703_846_fu_6863_p2;
wire   [15:0] add_ln703_847_fu_6868_p2;
wire   [15:0] add_ln703_866_fu_6972_p2;
wire   [15:0] sub_ln703_772_fu_6877_p2;
wire   [15:0] add_ln703_855_fu_6882_p2;
wire   [15:0] add_ln703_856_fu_6891_p2;
wire   [15:0] add_ln703_859_fu_6901_p2;
wire   [15:0] add_ln703_860_fu_6905_p2;
wire   [15:0] sub_ln703_775_fu_6910_p2;
wire   [15:0] add_ln703_861_fu_6919_p2;
wire   [15:0] add_ln703_862_fu_6923_p2;
wire   [15:0] sub_ln703_777_fu_6928_p2;
wire   [15:0] sub_ln703_778_fu_6933_p2;
wire   [15:0] sub_ln703_779_fu_6938_p2;
wire   [15:0] sub_ln703_782_fu_6946_p2;
wire   [15:0] sub_ln703_783_fu_6950_p2;
wire   [15:0] sub_ln703_784_fu_6954_p2;
wire   [15:0] sub_ln703_785_fu_6959_p2;
wire   [15:0] sub_ln703_786_fu_6964_p2;
wire   [15:0] add_ln703_865_fu_6968_p2;
wire   [15:0] add_ln703_869_fu_6976_p2;
wire   [15:0] sub_ln703_790_fu_6991_p2;
wire   [15:0] sub_ln703_791_fu_6996_p2;
wire   [15:0] sub_ln703_792_fu_7000_p2;
wire   [15:0] sub_ln703_793_fu_7005_p2;
wire   [15:0] sub_ln703_794_fu_7010_p2;
wire   [15:0] add_ln703_878_fu_7104_p2;
wire   [15:0] add_ln703_881_fu_7117_p2;
wire   [15:0] add_ln703_880_fu_7113_p2;
wire   [15:0] sub_ln703_795_fu_7015_p2;
wire   [15:0] sub_ln703_796_fu_7020_p2;
wire   [15:0] add_ln703_870_fu_7025_p2;
wire   [15:0] sub_ln703_798_fu_7035_p2;
wire   [15:0] sub_ln703_768_fu_6858_p2;
wire   [15:0] add_ln703_887_fu_7151_p2;
wire   [15:0] add_ln703_871_fu_7040_p2;
wire   [15:0] sub_ln703_800_fu_7045_p2;
wire   [15:0] sub_ln703_803_fu_7070_p2;
wire   [15:0] sub_ln703_804_fu_7075_p2;
wire   [15:0] sub_ln703_788_fu_6981_p2;
wire   [15:0] sub_ln703_773_fu_6886_p2;
wire   [15:0] sub_ln703_774_fu_6896_p2;
wire   [15:0] sub_ln703_806_fu_7089_p2;
wire   [15:0] add_ln703_879_fu_7108_p2;
wire   [15:0] add_ln703_883_fu_7127_p2;
wire   [15:0] add_ln703_885_fu_7142_p2;
wire   [15:0] add_ln703_886_fu_7147_p2;
wire   [15:0] add_ln703_889_fu_7161_p2;
wire   [15:0] sub_ln703_809_fu_7165_p2;
wire   [15:0] sub_ln703_810_fu_7170_p2;
wire   [15:0] sub_ln703_789_fu_6986_p2;
wire   [15:0] add_ln703_904_fu_7240_p2;
wire   [15:0] sub_ln703_780_fu_6942_p2;
wire   [15:0] add_ln703_909_fu_7255_p2;
wire   [15:0] add_ln703_908_fu_7250_p2;
wire   [15:0] add_ln703_916_fu_7269_p2;
wire   [15:0] add_ln703_915_fu_7265_p2;
wire   [15:0] add_ln703_921_fu_7283_p2;
wire   [15:0] add_ln703_919_fu_7279_p2;
wire   [15:0] sub_ln703_771_fu_6873_p2;
wire   [15:0] add_ln703_924_fu_7298_p2;
wire   [15:0] add_ln703_923_fu_7293_p2;
wire   [15:0] sub_ln703_776_fu_6915_p2;
wire   [15:0] add_ln703_931_fu_7308_p2;
wire   [15:0] add_ln703_910_fu_7259_p2;
wire   [15:0] add_ln703_925_fu_7302_p2;
wire   [15:0] add_ln703_932_fu_7313_p2;
wire   [15:0] sub_ln703_811_fu_7346_p2;
wire   [15:0] sub_ln703_812_fu_7350_p2;
wire   [15:0] add_ln703_890_fu_7354_p2;
wire   [15:0] add_ln703_891_fu_7358_p2;
wire   [15:0] add_ln703_897_fu_7362_p2;
wire   [15:0] add_ln703_899_fu_7366_p2;
wire   [15:0] sub_ln703_813_fu_7370_p2;
wire   [15:0] sub_ln703_815_fu_7374_p2;
wire   [15:0] add_ln703_900_fu_7378_p2;
wire   [15:0] add_ln703_901_fu_7390_p2;
wire   [15:0] add_ln703_902_fu_7394_p2;
wire   [15:0] sub_ln703_822_fu_7398_p2;
wire   [15:0] add_ln703_903_fu_7402_p2;
wire   [15:0] sub_ln703_826_fu_7407_p2;
wire   [15:0] sub_ln703_827_fu_7412_p2;
wire   [15:0] sub_ln703_828_fu_7417_p2;
wire   [15:0] sub_ln703_829_fu_7422_p2;
wire   [15:0] sub_ln703_831_fu_7430_p2;
wire   [15:0] sub_ln703_832_fu_7434_p2;
wire   [15:0] add_ln703_927_fu_7537_p2;
wire   [15:0] sub_ln703_833_fu_7439_p2;
wire   [15:0] sub_ln703_834_fu_7444_p2;
wire   [15:0] sub_ln703_836_fu_7453_p2;
wire   [15:0] sub_ln703_837_fu_7458_p2;
wire   [15:0] sub_ln703_839_fu_7467_p2;
wire   [15:0] add_ln703_907_fu_7477_p2;
wire   [15:0] add_ln703_911_fu_7481_p2;
wire   [15:0] sub_ln703_841_fu_7485_p2;
wire   [15:0] add_ln703_912_fu_7490_p2;
wire   [15:0] add_ln703_913_fu_7494_p2;
wire   [15:0] sub_ln703_842_fu_7498_p2;
wire   [15:0] sub_ln703_843_fu_7503_p2;
wire   [15:0] sub_ln703_844_fu_7508_p2;
wire   [15:0] add_ln703_918_fu_7513_p2;
wire   [15:0] sub_ln703_845_fu_7518_p2;
wire   [15:0] sub_ln703_846_fu_7523_p2;
wire   [15:0] sub_ln703_847_fu_7528_p2;
wire   [15:0] add_ln703_926_fu_7532_p2;
wire   [15:0] add_ln703_928_fu_7541_p2;
wire   [15:0] add_ln703_929_fu_7546_p2;
wire   [15:0] sub_ln703_848_fu_7551_p2;
wire   [15:0] add_ln703_937_fu_7659_p2;
wire   [15:0] sub_ln703_835_fu_7449_p2;
wire   [15:0] sub_ln703_849_fu_7556_p2;
wire   [15:0] add_ln703_930_fu_7561_p2;
wire   [15:0] sub_ln703_838_fu_7463_p2;
wire   [15:0] sub_ln703_850_fu_7566_p2;
wire   [15:0] sub_ln703_840_fu_7472_p2;
wire   [15:0] sub_ln703_851_fu_7571_p2;
wire   [15:0] sub_ln703_853_fu_7576_p2;
wire   [15:0] add_ln703_933_fu_7581_p2;
wire   [15:0] add_ln703_942_fu_7715_p2;
wire   [15:0] sub_ln703_855_fu_7591_p2;
wire   [15:0] sub_ln703_856_fu_7596_p2;
wire   [15:0] sub_ln703_860_fu_7620_p2;
wire   [15:0] sub_ln703_830_fu_7426_p2;
wire   [15:0] add_ln703_945_fu_7740_p2;
wire   [15:0] sub_ln703_861_fu_7625_p2;
wire   [15:0] add_ln703_935_fu_7629_p2;
wire   [15:0] sub_ln703_864_fu_7644_p2;
wire   [15:0] sub_ln703_817_fu_7382_p2;
wire   [15:0] add_ln703_950_fu_7770_p2;
wire   [15:0] add_ln703_949_fu_7765_p2;
wire   [15:0] add_ln703_940_fu_7690_p2;
wire   [15:0] sub_ln703_871_fu_7696_p2;
wire   [15:0] add_ln703_941_fu_7701_p2;
wire   [15:0] sub_ln703_872_fu_7705_p2;
wire   [15:0] sub_ln703_854_fu_7586_p2;
wire   [15:0] sub_ln703_874_fu_7725_p2;
wire   [15:0] add_ln703_947_fu_7745_p2;
wire   [15:0] add_ln703_957_fu_7823_p2;
wire   [15:0] add_ln703_956_fu_7819_p2;
wire   [15:0] add_ln703_951_fu_7774_p2;
wire   [15:0] add_ln703_952_fu_7800_p2;
wire   [15:0] add_ln703_955_fu_7815_p2;
wire   [15:0] sub_ln703_819_fu_7386_p2;
wire   [15:0] add_ln703_1000_fu_7852_p2;
wire   [15:0] add_ln703_1002_fu_7863_p2;
wire   [15:0] add_ln703_1003_fu_7867_p2;
wire   [15:0] add_ln703_1001_fu_7857_p2;
wire   [15:0] sub_ln703_876_fu_7878_p2;
wire   [15:0] add_ln703_944_fu_7882_p2;
wire   [15:0] sub_ln703_877_fu_7886_p2;
wire   [15:0] sub_ln703_878_fu_7890_p2;
wire   [15:0] sub_ln703_883_fu_7898_p2;
wire   [15:0] sub_ln703_885_fu_7906_p2;
wire   [15:0] sub_ln703_888_fu_7918_p2;
wire   [15:0] sub_ln703_889_fu_7922_p2;
wire   [15:0] sub_ln703_890_fu_7926_p2;
wire   [15:0] sub_ln703_891_fu_7930_p2;
wire   [15:0] sub_ln703_896_fu_7934_p2;
wire   [15:0] add_ln703_953_fu_7956_p2;
wire   [15:0] sub_ln703_902_fu_7961_p2;
wire   [15:0] sub_ln703_903_fu_7966_p2;
wire   [15:0] sub_ln703_905_fu_7970_p2;
wire   [15:0] sub_ln703_906_fu_7974_p2;
wire   [15:0] sub_ln703_908_fu_7983_p2;
wire   [15:0] sub_ln703_886_fu_7910_p2;
wire   [15:0] add_ln703_959_fu_7997_p2;
wire   [15:0] sub_ln703_913_fu_8007_p2;
wire   [15:0] add_ln703_960_fu_8012_p2;
wire   [15:0] add_ln703_961_fu_8016_p2;
wire   [15:0] sub_ln703_914_fu_8020_p2;
wire   [15:0] sub_ln703_915_fu_8024_p2;
wire   [15:0] sub_ln703_897_fu_7938_p2;
wire   [15:0] sub_ln703_918_fu_8033_p2;
wire   [15:0] sub_ln703_921_fu_8047_p2;
wire   [15:0] add_ln703_970_fu_8125_p2;
wire   [15:0] add_ln703_962_fu_8052_p2;
wire   [15:0] sub_ln703_923_fu_8057_p2;
wire   [15:0] sub_ln703_882_fu_7894_p2;
wire   [15:0] add_ln703_972_fu_8148_p2;
wire   [15:0] sub_ln703_907_fu_7978_p2;
wire   [15:0] add_ln703_963_fu_8062_p2;
wire   [15:0] sub_ln703_884_fu_7902_p2;
wire   [15:0] add_ln703_975_fu_8170_p2;
wire   [15:0] add_ln703_965_fu_8067_p2;
wire   [15:0] sub_ln703_887_fu_7914_p2;
wire   [15:0] add_ln703_977_fu_8186_p2;
wire   [15:0] sub_ln703_910_fu_7992_p2;
wire   [15:0] sub_ln703_912_fu_8002_p2;
wire   [15:0] sub_ln703_928_fu_8090_p2;
wire   [15:0] sub_ln703_929_fu_8095_p2;
wire   [15:0] add_ln703_966_fu_8100_p2;
wire   [15:0] add_ln703_967_fu_8105_p2;
wire   [15:0] add_ln703_968_fu_8110_p2;
wire   [15:0] add_ln703_969_fu_8115_p2;
wire   [15:0] sub_ln703_899_fu_7942_p2;
wire   [15:0] add_ln703_982_fu_8239_p2;
wire   [15:0] sub_ln703_900_fu_7946_p2;
wire   [15:0] add_ln703_984_fu_8250_p2;
wire   [15:0] sub_ln703_901_fu_7951_p2;
wire   [15:0] add_ln703_987_fu_8260_p2;
wire   [15:0] sub_ln703_919_fu_8037_p2;
wire   [15:0] sub_ln703_920_fu_8042_p2;
wire   [15:0] sub_ln703_930_fu_8120_p2;
wire   [15:0] add_ln703_971_fu_8129_p2;
wire   [15:0] sub_ln703_931_fu_8134_p2;
wire   [15:0] sub_ln703_932_fu_8139_p2;
wire   [15:0] sub_ln703_933_fu_8143_p2;
wire   [15:0] add_ln703_973_fu_8153_p2;
wire   [15:0] add_ln703_974_fu_8159_p2;
wire   [15:0] sub_ln703_934_fu_8165_p2;
wire   [15:0] add_ln703_976_fu_8175_p2;
wire   [15:0] sub_ln703_909_fu_7987_p2;
wire   [15:0] add_ln703_994_fu_8325_p2;
wire   [15:0] sub_ln703_935_fu_8181_p2;
wire   [15:0] add_ln703_978_fu_8191_p2;
wire   [15:0] add_ln703_979_fu_8197_p2;
wire   [15:0] sub_ln703_924_fu_8072_p2;
wire   [15:0] sub_ln703_925_fu_8076_p2;
wire   [15:0] sub_ln703_926_fu_8080_p2;
wire   [15:0] add_ln703_980_fu_8203_p2;
wire   [15:0] sub_ln703_927_fu_8085_p2;
wire   [15:0] sub_ln703_936_fu_8209_p2;
wire   [15:0] add_ln703_981_fu_8214_p2;
wire   [15:0] sub_ln703_937_fu_8219_p2;
wire   [15:0] sub_ln703_938_fu_8224_p2;
wire   [15:0] sub_ln703_916_fu_8028_p2;
wire   [15:0] add_ln703_1007_fu_8395_p2;
wire   [15:0] sub_ln703_939_fu_8229_p2;
wire   [15:0] add_ln703_1009_fu_8410_p2;
wire   [15:0] sub_ln703_940_fu_8234_p2;
wire   [15:0] add_ln703_983_fu_8244_p2;
wire   [15:0] add_ln703_986_fu_8255_p2;
wire   [15:0] acc_1_V_fu_8265_p2;
wire   [15:0] acc_2_V_fu_8270_p2;
wire   [15:0] acc_3_V_fu_8275_p2;
wire   [15:0] acc_4_V_fu_8280_p2;
wire   [15:0] acc_5_V_fu_8285_p2;
wire   [15:0] acc_6_V_fu_8290_p2;
wire   [15:0] acc_7_V_fu_8295_p2;
wire   [15:0] acc_8_V_fu_8300_p2;
wire   [15:0] acc_9_V_fu_8305_p2;
wire   [15:0] acc_10_V_fu_8310_p2;
wire   [15:0] acc_11_V_fu_8315_p2;
wire   [15:0] acc_12_V_fu_8320_p2;
wire   [15:0] acc_13_V_fu_8330_p2;
wire   [15:0] acc_14_V_fu_8335_p2;
wire   [15:0] acc_15_V_fu_8340_p2;
wire   [15:0] acc_16_V_fu_8345_p2;
wire   [15:0] acc_17_V_fu_8350_p2;
wire   [15:0] acc_18_V_fu_8355_p2;
wire   [15:0] acc_19_V_fu_8360_p2;
wire   [15:0] acc_20_V_fu_8365_p2;
wire   [15:0] acc_22_V_fu_8370_p2;
wire   [15:0] acc_23_V_fu_8375_p2;
wire   [15:0] acc_24_V_fu_8380_p2;
wire   [15:0] acc_25_V_fu_8385_p2;
wire   [15:0] acc_26_V_fu_8390_p2;
wire   [15:0] acc_27_V_fu_8400_p2;
wire   [15:0] acc_28_V_fu_8405_p2;
wire   [15:0] acc_29_V_fu_8414_p2;
wire   [15:0] acc_30_V_fu_8419_p2;
wire   [15:0] acc_31_V_fu_8424_p2;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] data_32_V_read_int_reg;
reg   [15:0] data_33_V_read_int_reg;
reg   [15:0] data_34_V_read_int_reg;
reg   [15:0] data_35_V_read_int_reg;
reg   [15:0] data_36_V_read_int_reg;
reg   [15:0] data_37_V_read_int_reg;
reg   [15:0] data_38_V_read_int_reg;
reg   [15:0] data_39_V_read_int_reg;
reg   [15:0] data_40_V_read_int_reg;
reg   [15:0] data_41_V_read_int_reg;
reg   [15:0] data_42_V_read_int_reg;
reg   [15:0] data_43_V_read_int_reg;
reg   [15:0] data_44_V_read_int_reg;
reg   [15:0] data_45_V_read_int_reg;
reg   [15:0] data_46_V_read_int_reg;
reg   [15:0] data_47_V_read_int_reg;
reg   [15:0] data_48_V_read_int_reg;
reg   [15:0] data_49_V_read_int_reg;
reg   [15:0] data_50_V_read_int_reg;
reg   [15:0] data_51_V_read_int_reg;
reg   [15:0] data_52_V_read_int_reg;
reg   [15:0] data_53_V_read_int_reg;
reg   [15:0] data_54_V_read_int_reg;
reg   [15:0] data_55_V_read_int_reg;
reg   [15:0] data_56_V_read_int_reg;
reg   [15:0] data_57_V_read_int_reg;
reg   [15:0] data_58_V_read_int_reg;
reg   [15:0] data_59_V_read_int_reg;
reg   [15:0] data_60_V_read_int_reg;
reg   [15:0] data_61_V_read_int_reg;
reg   [15:0] data_62_V_read_int_reg;
reg   [15:0] data_63_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        acc_21_V_reg_12991 <= acc_21_V_fu_7872_p2;
        add_ln703_130_reg_10373 <= add_ln703_130_fu_556_p2;
        add_ln703_131_reg_10354 <= add_ln703_131_fu_544_p2;
        add_ln703_131_reg_10354_pp0_iter2_reg <= add_ln703_131_reg_10354;
        add_ln703_132_reg_10414 <= add_ln703_132_fu_599_p2;
        add_ln703_134_reg_10385 <= add_ln703_134_fu_568_p2;
        add_ln703_135_reg_10425 <= add_ln703_135_fu_619_p2;
        add_ln703_140_reg_10442 <= add_ln703_140_fu_644_p2;
        add_ln703_141_reg_10447 <= add_ln703_141_fu_649_p2;
        add_ln703_144_reg_10403 <= add_ln703_144_fu_589_p2;
        add_ln703_144_reg_10403_pp0_iter3_reg <= add_ln703_144_reg_10403;
        add_ln703_153_reg_10503 <= add_ln703_153_fu_809_p2;
        add_ln703_157_reg_10529 <= add_ln703_157_fu_892_p2;
        add_ln703_158_reg_10482 <= add_ln703_158_fu_676_p2;
        add_ln703_161_reg_10487 <= add_ln703_161_fu_681_p2;
        add_ln703_162_reg_10539 <= add_ln703_162_fu_917_p2;
        add_ln703_170_reg_10566 <= add_ln703_170_fu_972_p2;
        add_ln703_171_reg_10571 <= add_ln703_171_fu_977_p2;
        add_ln703_173_reg_10576 <= add_ln703_173_fu_982_p2;
        add_ln703_177_reg_10591 <= add_ln703_177_fu_997_p2;
        add_ln703_179_reg_10495 <= add_ln703_179_fu_685_p2;
        add_ln703_181_reg_10601 <= add_ln703_181_fu_1015_p2;
        add_ln703_183_reg_10606 <= add_ln703_183_fu_1021_p2;
        add_ln703_186_reg_10621 <= add_ln703_186_fu_1036_p2;
        add_ln703_192_reg_10626 <= add_ln703_192_fu_1050_p2;
        add_ln703_204_reg_10641 <= add_ln703_204_fu_1059_p2;
        add_ln703_207_reg_10682 <= add_ln703_207_fu_1299_p2;
        add_ln703_208_reg_10687 <= add_ln703_208_fu_1309_p2;
        add_ln703_209_reg_10646 <= add_ln703_209_fu_1064_p2;
        add_ln703_210_reg_10692 <= add_ln703_210_fu_1314_p2;
        add_ln703_213_reg_10653 <= add_ln703_213_fu_1068_p2;
        add_ln703_216_reg_10702 <= add_ln703_216_fu_1358_p2;
        add_ln703_223_reg_10658 <= add_ln703_223_fu_1073_p2;
        add_ln703_224_reg_10732 <= add_ln703_224_fu_1437_p2;
        add_ln703_226_reg_10737 <= add_ln703_226_fu_1457_p2;
        add_ln703_227_reg_10752 <= add_ln703_227_fu_1472_p2;
        add_ln703_233_reg_10767 <= add_ln703_233_fu_1501_p2;
        add_ln703_236_reg_10772 <= add_ln703_236_fu_1511_p2;
        add_ln703_238_reg_10777 <= add_ln703_238_fu_1520_p2;
        add_ln703_247_reg_10802 <= add_ln703_247_fu_1563_p2;
        add_ln703_250_reg_10807 <= add_ln703_250_fu_1574_p2;
        add_ln703_252_reg_10665 <= add_ln703_252_fu_1077_p2;
        add_ln703_252_reg_10665_pp0_iter5_reg <= add_ln703_252_reg_10665;
        add_ln703_254_reg_10672 <= add_ln703_254_fu_1081_p2;
        add_ln703_260_reg_10817 <= add_ln703_260_fu_1593_p2;
        add_ln703_262_reg_10827 <= add_ln703_262_fu_1604_p2;
        add_ln703_265_reg_10837 <= add_ln703_265_fu_1614_p2;
        add_ln703_280_reg_10846 <= add_ln703_280_fu_1618_p2;
        add_ln703_283_reg_10873 <= add_ln703_283_fu_1979_p2;
        add_ln703_285_reg_10888 <= add_ln703_285_fu_2009_p2;
        add_ln703_289_reg_10898 <= add_ln703_289_fu_2034_p2;
        add_ln703_290_reg_10903 <= add_ln703_290_fu_2039_p2;
        add_ln703_294_reg_10918 <= add_ln703_294_fu_2084_p2;
        add_ln703_295_reg_10923 <= add_ln703_295_fu_2089_p2;
        add_ln703_300_reg_10930 <= add_ln703_300_fu_2093_p2;
        add_ln703_303_reg_10940 <= add_ln703_303_fu_2104_p2;
        add_ln703_304_reg_10945 <= add_ln703_304_fu_2110_p2;
        add_ln703_307_reg_10960 <= add_ln703_307_fu_2125_p2;
        add_ln703_309_reg_10970 <= add_ln703_309_fu_2136_p2;
        add_ln703_310_reg_10980 <= add_ln703_310_fu_2147_p2;
        add_ln703_323_reg_11005 <= add_ln703_323_fu_2188_p2;
        add_ln703_326_reg_10855 <= add_ln703_326_fu_1622_p2;
        add_ln703_326_reg_10855_pp0_iter6_reg <= add_ln703_326_reg_10855;
        add_ln703_328_reg_11015 <= add_ln703_328_fu_2208_p2;
        add_ln703_333_reg_11025 <= add_ln703_333_fu_2224_p2;
        add_ln703_341_reg_11030 <= add_ln703_341_fu_2230_p2;
        add_ln703_342_reg_11071 <= add_ln703_342_fu_2520_p2;
        add_ln703_346_reg_11106 <= add_ln703_346_fu_2589_p2;
        add_ln703_350_reg_11111 <= add_ln703_350_fu_2602_p2;
        add_ln703_352_reg_11126 <= add_ln703_352_fu_2633_p2;
        add_ln703_354_reg_11131 <= add_ln703_354_fu_2638_p2;
        add_ln703_356_reg_11148 <= add_ln703_356_fu_2657_p2;
        add_ln703_360_reg_11158 <= add_ln703_360_fu_2677_p2;
        add_ln703_369_reg_11037 <= add_ln703_369_fu_2234_p2;
        add_ln703_369_reg_11037_pp0_iter7_reg <= add_ln703_369_reg_11037;
        add_ln703_371_reg_11193 <= add_ln703_371_fu_2732_p2;
        add_ln703_375_reg_11198 <= add_ln703_375_fu_2738_p2;
        add_ln703_384_reg_11203 <= add_ln703_384_fu_2743_p2;
        add_ln703_386_reg_11262 <= add_ln703_386_fu_3015_p2;
        add_ln703_390_reg_11272 <= add_ln703_390_fu_3050_p2;
        add_ln703_400_reg_11210 <= add_ln703_400_fu_2752_p2;
        add_ln703_402_reg_11215 <= add_ln703_402_fu_2758_p2;
        add_ln703_402_reg_11215_pp0_iter8_reg <= add_ln703_402_reg_11215;
        add_ln703_410_reg_11287 <= add_ln703_410_fu_3149_p2;
        add_ln703_416_reg_11297 <= add_ln703_416_fu_3170_p2;
        add_ln703_417_reg_11312 <= add_ln703_417_fu_3185_p2;
        add_ln703_424_reg_11225 <= add_ln703_424_fu_2762_p2;
        add_ln703_426_reg_11347 <= add_ln703_426_fu_3258_p2;
        add_ln703_431_reg_11357 <= add_ln703_431_fu_3274_p2;
        add_ln703_435_reg_11362 <= add_ln703_435_fu_3284_p2;
        add_ln703_438_reg_11382 <= add_ln703_438_fu_3310_p2;
        add_ln703_439_reg_11233 <= add_ln703_439_fu_2766_p2;
        add_ln703_439_reg_11233_pp0_iter8_reg <= add_ln703_439_reg_11233;
        add_ln703_445_reg_11387 <= add_ln703_445_fu_3315_p2;
        add_ln703_447_reg_11392 <= add_ln703_447_fu_3320_p2;
        add_ln703_451_reg_11402 <= add_ln703_451_fu_3329_p2;
        add_ln703_466_reg_11410 <= add_ln703_466_fu_3333_p2;
        add_ln703_469_reg_11479 <= add_ln703_469_fu_3655_p2;
        add_ln703_471_reg_11418 <= add_ln703_471_fu_3337_p2;
        add_ln703_476_reg_11494 <= add_ln703_476_fu_3685_p2;
        add_ln703_478_reg_11519 <= add_ln703_478_fu_3730_p2;
        add_ln703_484_reg_11423 <= add_ln703_484_fu_3342_p2;
        add_ln703_490_reg_11428 <= add_ln703_490_fu_3347_p2;
        add_ln703_496_reg_11544 <= add_ln703_496_fu_3806_p2;
        add_ln703_497_reg_11549 <= add_ln703_497_fu_3811_p2;
        add_ln703_498_reg_11436 <= add_ln703_498_fu_3351_p2;
        add_ln703_506_reg_11559 <= add_ln703_506_fu_3839_p2;
        add_ln703_507_reg_11441 <= add_ln703_507_fu_3356_p2;
        add_ln703_507_reg_11441_pp0_iter9_reg <= add_ln703_507_reg_11441;
        add_ln703_512_reg_11589 <= add_ln703_512_fu_3878_p2;
        add_ln703_515_reg_11599 <= add_ln703_515_fu_3889_p2;
        add_ln703_517_reg_11604 <= add_ln703_517_fu_3894_p2;
        add_ln703_525_reg_11243 <= add_ln703_525_fu_2774_p2;
        add_ln703_525_reg_11243_pp0_iter8_reg <= add_ln703_525_reg_11243;
        add_ln703_525_reg_11243_pp0_iter9_reg <= add_ln703_525_reg_11243_pp0_iter8_reg;
        add_ln703_528_reg_11452 <= add_ln703_528_fu_3360_p2;
        add_ln703_528_reg_11452_pp0_iter9_reg <= add_ln703_528_reg_11452;
        add_ln703_534_reg_11248 <= add_ln703_534_fu_2779_p2;
        add_ln703_534_reg_11248_pp0_iter8_reg <= add_ln703_534_reg_11248;
        add_ln703_534_reg_11248_pp0_iter9_reg <= add_ln703_534_reg_11248_pp0_iter8_reg;
        add_ln703_535_reg_11457 <= add_ln703_535_fu_3364_p2;
        add_ln703_537_reg_11609 <= add_ln703_537_fu_3912_p2;
        add_ln703_545_reg_11614 <= add_ln703_545_fu_3923_p2;
        add_ln703_556_reg_11619 <= add_ln703_556_fu_3933_p2;
        add_ln703_560_reg_11629 <= add_ln703_560_fu_3943_p2;
        add_ln703_566_reg_11635 <= add_ln703_566_fu_3952_p2;
        add_ln703_568_reg_11464 <= add_ln703_568_fu_3368_p2;
        add_ln703_568_reg_11464_pp0_iter9_reg <= add_ln703_568_reg_11464;
        add_ln703_569_reg_11640 <= add_ln703_569_fu_3957_p2;
        add_ln703_572_reg_11698 <= add_ln703_572_fu_4308_p2;
        add_ln703_573_reg_11708 <= add_ln703_573_fu_4323_p2;
        add_ln703_581_reg_11723 <= add_ln703_581_fu_4358_p2;
        add_ln703_583_reg_11728 <= add_ln703_583_fu_4363_p2;
        add_ln703_586_reg_11743 <= add_ln703_586_fu_4398_p2;
        add_ln703_588_reg_11646 <= add_ln703_588_fu_3961_p2;
        add_ln703_590_reg_11748 <= add_ln703_590_fu_4412_p2;
        add_ln703_591_reg_11758 <= add_ln703_591_fu_4423_p2;
        add_ln703_592_reg_11763 <= add_ln703_592_fu_4428_p2;
        add_ln703_598_reg_11768 <= add_ln703_598_fu_4441_p2;
        add_ln703_599_reg_11798 <= add_ln703_599_fu_4477_p2;
        add_ln703_600_reg_11652 <= add_ln703_600_fu_3965_p2;
        add_ln703_600_reg_11652_pp0_iter10_reg <= add_ln703_600_reg_11652;
        add_ln703_609_reg_11803 <= add_ln703_609_fu_4501_p2;
        add_ln703_616_reg_11808 <= add_ln703_616_fu_4511_p2;
        add_ln703_621_reg_11662 <= add_ln703_621_fu_3969_p2;
        add_ln703_621_reg_11662_pp0_iter10_reg <= add_ln703_621_reg_11662;
        add_ln703_633_reg_11823 <= add_ln703_633_fu_4531_p2;
        add_ln703_634_reg_11828 <= add_ln703_634_fu_4535_p2;
        add_ln703_639_reg_11833 <= add_ln703_639_fu_4541_p2;
        add_ln703_646_reg_11838 <= add_ln703_646_fu_4546_p2;
        add_ln703_647_reg_11874 <= add_ln703_647_fu_4870_p2;
        add_ln703_648_reg_11889 <= add_ln703_648_fu_4899_p2;
        add_ln703_650_reg_11844 <= add_ln703_650_fu_4550_p2;
        add_ln703_650_reg_11844_pp0_iter11_reg <= add_ln703_650_reg_11844;
        add_ln703_651_reg_11929 <= add_ln703_651_fu_4959_p2;
        add_ln703_660_reg_11939 <= add_ln703_660_fu_4994_p2;
        add_ln703_661_reg_11944 <= add_ln703_661_fu_4999_p2;
        add_ln703_666_reg_11954 <= add_ln703_666_fu_5013_p2;
        add_ln703_667_reg_11853 <= add_ln703_667_fu_4554_p2;
        add_ln703_668_reg_11959 <= add_ln703_668_fu_5019_p2;
        add_ln703_676_reg_11979 <= add_ln703_676_fu_5052_p2;
        add_ln703_682_reg_11984 <= add_ln703_682_fu_5066_p2;
        add_ln703_685_reg_11989 <= add_ln703_685_fu_5077_p2;
        add_ln703_691_reg_11994 <= add_ln703_691_fu_5092_p2;
        add_ln703_697_reg_12002 <= add_ln703_697_fu_5096_p2;
        add_ln703_703_reg_12022 <= add_ln703_703_fu_5116_p2;
        add_ln703_704_reg_12056 <= add_ln703_704_fu_5336_p2;
        add_ln703_706_reg_12031 <= add_ln703_706_fu_5120_p2;
        add_ln703_719_reg_12086 <= add_ln703_719_fu_5439_p2;
        add_ln703_722_reg_12036 <= add_ln703_722_fu_5125_p2;
        add_ln703_726_reg_12041 <= add_ln703_726_fu_5130_p2;
        add_ln703_728_reg_12096 <= add_ln703_728_fu_5485_p2;
        add_ln703_733_reg_12146 <= add_ln703_733_fu_5551_p2;
        add_ln703_734_reg_12151 <= add_ln703_734_fu_5556_p2;
        add_ln703_735_reg_12161 <= add_ln703_735_fu_5571_p2;
        add_ln703_737_reg_12047 <= add_ln703_737_fu_5134_p2;
        add_ln703_755_reg_12196 <= add_ln703_755_fu_5652_p2;
        add_ln703_765_reg_12219 <= add_ln703_765_fu_5671_p2;
        add_ln703_770_reg_12258 <= add_ln703_770_fu_5950_p2;
        add_ln703_778_reg_12227 <= add_ln703_778_fu_5675_p2;
        add_ln703_779_reg_12273 <= add_ln703_779_fu_6024_p2;
        add_ln703_783_reg_12236 <= add_ln703_783_fu_5679_p2;
        add_ln703_791_reg_12348 <= add_ln703_791_fu_6131_p2;
        add_ln703_792_reg_12363 <= add_ln703_792_fu_6146_p2;
        add_ln703_796_reg_12368 <= add_ln703_796_fu_6160_p2;
        add_ln703_798_reg_12373 <= add_ln703_798_fu_6166_p2;
        add_ln703_801_reg_12393 <= add_ln703_801_fu_6187_p2;
        add_ln703_802_reg_12398 <= add_ln703_802_fu_6192_p2;
        add_ln703_816_reg_12241 <= add_ln703_816_fu_5684_p2;
        add_ln703_816_reg_12241_pp0_iter13_reg <= add_ln703_816_reg_12241;
        add_ln703_818_reg_12409 <= add_ln703_818_fu_6205_p2;
        add_ln703_818_reg_12409_pp0_iter14_reg <= add_ln703_818_reg_12409;
        add_ln703_819_reg_12455 <= add_ln703_819_fu_6447_p2;
        add_ln703_821_reg_12414 <= add_ln703_821_fu_6216_p2;
        add_ln703_825_reg_12480 <= add_ln703_825_fu_6526_p2;
        add_ln703_826_reg_12419 <= add_ln703_826_fu_6222_p2;
        add_ln703_827_reg_12485 <= add_ln703_827_fu_6531_p2;
        add_ln703_831_reg_12490 <= add_ln703_831_fu_6554_p2;
        add_ln703_833_reg_12495 <= add_ln703_833_fu_6573_p2;
        add_ln703_834_reg_12505 <= add_ln703_834_fu_6594_p2;
        add_ln703_836_reg_12428 <= add_ln703_836_fu_6226_p2;
        add_ln703_838_reg_12520 <= add_ln703_838_fu_6634_p2;
        add_ln703_840_reg_12535 <= add_ln703_840_fu_6649_p2;
        add_ln703_841_reg_12550 <= add_ln703_841_fu_6664_p2;
        add_ln703_845_reg_12560 <= add_ln703_845_fu_6689_p2;
        add_ln703_849_reg_12434 <= add_ln703_849_fu_6230_p2;
        add_ln703_849_reg_12434_pp0_iter14_reg <= add_ln703_849_reg_12434;
        add_ln703_851_reg_12565 <= add_ln703_851_fu_6702_p2;
        add_ln703_858_reg_12575 <= add_ln703_858_fu_6733_p2;
        add_ln703_867_reg_12444 <= add_ln703_867_fu_6234_p2;
        add_ln703_867_reg_12444_pp0_iter14_reg <= add_ln703_867_reg_12444;
        add_ln703_868_reg_12585 <= add_ln703_868_fu_6755_p2;
        add_ln703_872_reg_12650 <= add_ln703_872_fu_7050_p2;
        add_ln703_873_reg_12655 <= add_ln703_873_fu_7055_p2;
        add_ln703_874_reg_12675 <= add_ln703_874_fu_7084_p2;
        add_ln703_875_reg_12680 <= add_ln703_875_fu_7094_p2;
        add_ln703_876_reg_12600 <= add_ln703_876_fu_6769_p2;
        add_ln703_877_reg_12605 <= add_ln703_877_fu_6774_p2;
        add_ln703_882_reg_12690 <= add_ln703_882_fu_7121_p2;
        add_ln703_884_reg_12695 <= add_ln703_884_fu_7132_p2;
        add_ln703_888_reg_12705 <= add_ln703_888_fu_7156_p2;
        add_ln703_892_reg_12710 <= add_ln703_892_fu_7175_p2;
        add_ln703_893_reg_12715 <= add_ln703_893_fu_7180_p2;
        add_ln703_894_reg_12616 <= add_ln703_894_fu_6778_p2;
        add_ln703_894_reg_12616_pp0_iter15_reg <= add_ln703_894_reg_12616;
        add_ln703_895_reg_12720 <= add_ln703_895_fu_7185_p2;
        add_ln703_896_reg_12725 <= add_ln703_896_fu_7190_p2;
        add_ln703_898_reg_12730 <= add_ln703_898_fu_7195_p2;
        add_ln703_905_reg_12625 <= add_ln703_905_fu_6782_p2;
        add_ln703_906_reg_12775 <= add_ln703_906_fu_7245_p2;
        add_ln703_914_reg_12632 <= add_ln703_914_fu_6786_p2;
        add_ln703_917_reg_12780 <= add_ln703_917_fu_7273_p2;
        add_ln703_920_reg_12637 <= add_ln703_920_fu_6791_p2;
        add_ln703_920_reg_12637_pp0_iter15_reg <= add_ln703_920_reg_12637;
        add_ln703_922_reg_12785 <= add_ln703_922_fu_7287_p2;
        add_ln703_934_reg_12845 <= add_ln703_934_fu_7610_p2;
        add_ln703_936_reg_12855 <= add_ln703_936_fu_7634_p2;
        add_ln703_938_reg_12875 <= add_ln703_938_fu_7663_p2;
        add_ln703_939_reg_12890 <= add_ln703_939_fu_7679_p2;
        add_ln703_943_reg_12905 <= add_ln703_943_fu_7719_p2;
        add_ln703_946_reg_12805 <= add_ln703_946_fu_7334_p2;
        add_ln703_948_reg_12930 <= add_ln703_948_fu_7760_p2;
        add_ln703_954_reg_12812 <= add_ln703_954_fu_7338_p2;
        add_ln703_958_reg_12965 <= add_ln703_958_fu_7827_p2;
        add_ln703_964_reg_12985 <= add_ln703_964_fu_7848_p2;
        add_ln703_985_reg_12819 <= add_ln703_985_fu_7342_p2;
        add_ln703_985_reg_12819_pp0_iter16_reg <= add_ln703_985_reg_12819;
        add_ln703_reg_10335 <= add_ln703_fu_530_p2;
        add_ln703_reg_10335_pp0_iter1_reg <= add_ln703_reg_10335;
        data_0_V_read_10_reg_10329 <= data_0_V_read_int_reg;
        data_10_V_read11_reg_10105 <= data_10_V_read_int_reg;
        data_10_V_read11_reg_10105_pp0_iter1_reg <= data_10_V_read11_reg_10105;
        data_10_V_read11_reg_10105_pp0_iter2_reg <= data_10_V_read11_reg_10105_pp0_iter1_reg;
        data_10_V_read11_reg_10105_pp0_iter3_reg <= data_10_V_read11_reg_10105_pp0_iter2_reg;
        data_10_V_read11_reg_10105_pp0_iter4_reg <= data_10_V_read11_reg_10105_pp0_iter3_reg;
        data_11_V_read12_reg_10075 <= data_11_V_read_int_reg;
        data_11_V_read12_reg_10075_pp0_iter1_reg <= data_11_V_read12_reg_10075;
        data_11_V_read12_reg_10075_pp0_iter2_reg <= data_11_V_read12_reg_10075_pp0_iter1_reg;
        data_11_V_read12_reg_10075_pp0_iter3_reg <= data_11_V_read12_reg_10075_pp0_iter2_reg;
        data_11_V_read12_reg_10075_pp0_iter4_reg <= data_11_V_read12_reg_10075_pp0_iter3_reg;
        data_11_V_read12_reg_10075_pp0_iter5_reg <= data_11_V_read12_reg_10075_pp0_iter4_reg;
        data_12_V_read13_reg_10045 <= data_12_V_read_int_reg;
        data_12_V_read13_reg_10045_pp0_iter1_reg <= data_12_V_read13_reg_10045;
        data_12_V_read13_reg_10045_pp0_iter2_reg <= data_12_V_read13_reg_10045_pp0_iter1_reg;
        data_12_V_read13_reg_10045_pp0_iter3_reg <= data_12_V_read13_reg_10045_pp0_iter2_reg;
        data_12_V_read13_reg_10045_pp0_iter4_reg <= data_12_V_read13_reg_10045_pp0_iter3_reg;
        data_12_V_read13_reg_10045_pp0_iter5_reg <= data_12_V_read13_reg_10045_pp0_iter4_reg;
        data_13_V_read14_reg_10015 <= data_13_V_read_int_reg;
        data_13_V_read14_reg_10015_pp0_iter1_reg <= data_13_V_read14_reg_10015;
        data_13_V_read14_reg_10015_pp0_iter2_reg <= data_13_V_read14_reg_10015_pp0_iter1_reg;
        data_13_V_read14_reg_10015_pp0_iter3_reg <= data_13_V_read14_reg_10015_pp0_iter2_reg;
        data_13_V_read14_reg_10015_pp0_iter4_reg <= data_13_V_read14_reg_10015_pp0_iter3_reg;
        data_13_V_read14_reg_10015_pp0_iter5_reg <= data_13_V_read14_reg_10015_pp0_iter4_reg;
        data_14_V_read15_reg_9987 <= data_14_V_read_int_reg;
        data_14_V_read15_reg_9987_pp0_iter1_reg <= data_14_V_read15_reg_9987;
        data_14_V_read15_reg_9987_pp0_iter2_reg <= data_14_V_read15_reg_9987_pp0_iter1_reg;
        data_14_V_read15_reg_9987_pp0_iter3_reg <= data_14_V_read15_reg_9987_pp0_iter2_reg;
        data_14_V_read15_reg_9987_pp0_iter4_reg <= data_14_V_read15_reg_9987_pp0_iter3_reg;
        data_14_V_read15_reg_9987_pp0_iter5_reg <= data_14_V_read15_reg_9987_pp0_iter4_reg;
        data_15_V_read16_reg_9962 <= data_15_V_read_int_reg;
        data_15_V_read16_reg_9962_pp0_iter1_reg <= data_15_V_read16_reg_9962;
        data_15_V_read16_reg_9962_pp0_iter2_reg <= data_15_V_read16_reg_9962_pp0_iter1_reg;
        data_15_V_read16_reg_9962_pp0_iter3_reg <= data_15_V_read16_reg_9962_pp0_iter2_reg;
        data_15_V_read16_reg_9962_pp0_iter4_reg <= data_15_V_read16_reg_9962_pp0_iter3_reg;
        data_15_V_read16_reg_9962_pp0_iter5_reg <= data_15_V_read16_reg_9962_pp0_iter4_reg;
        data_16_V_read17_reg_9935 <= data_16_V_read_int_reg;
        data_16_V_read17_reg_9935_pp0_iter1_reg <= data_16_V_read17_reg_9935;
        data_16_V_read17_reg_9935_pp0_iter2_reg <= data_16_V_read17_reg_9935_pp0_iter1_reg;
        data_16_V_read17_reg_9935_pp0_iter3_reg <= data_16_V_read17_reg_9935_pp0_iter2_reg;
        data_16_V_read17_reg_9935_pp0_iter4_reg <= data_16_V_read17_reg_9935_pp0_iter3_reg;
        data_16_V_read17_reg_9935_pp0_iter5_reg <= data_16_V_read17_reg_9935_pp0_iter4_reg;
        data_16_V_read17_reg_9935_pp0_iter6_reg <= data_16_V_read17_reg_9935_pp0_iter5_reg;
        data_17_V_read18_reg_9904 <= data_17_V_read_int_reg;
        data_17_V_read18_reg_9904_pp0_iter1_reg <= data_17_V_read18_reg_9904;
        data_17_V_read18_reg_9904_pp0_iter2_reg <= data_17_V_read18_reg_9904_pp0_iter1_reg;
        data_17_V_read18_reg_9904_pp0_iter3_reg <= data_17_V_read18_reg_9904_pp0_iter2_reg;
        data_17_V_read18_reg_9904_pp0_iter4_reg <= data_17_V_read18_reg_9904_pp0_iter3_reg;
        data_17_V_read18_reg_9904_pp0_iter5_reg <= data_17_V_read18_reg_9904_pp0_iter4_reg;
        data_17_V_read18_reg_9904_pp0_iter6_reg <= data_17_V_read18_reg_9904_pp0_iter5_reg;
        data_18_V_read_8_reg_9874 <= data_18_V_read_int_reg;
        data_18_V_read_8_reg_9874_pp0_iter1_reg <= data_18_V_read_8_reg_9874;
        data_18_V_read_8_reg_9874_pp0_iter2_reg <= data_18_V_read_8_reg_9874_pp0_iter1_reg;
        data_18_V_read_8_reg_9874_pp0_iter3_reg <= data_18_V_read_8_reg_9874_pp0_iter2_reg;
        data_18_V_read_8_reg_9874_pp0_iter4_reg <= data_18_V_read_8_reg_9874_pp0_iter3_reg;
        data_18_V_read_8_reg_9874_pp0_iter5_reg <= data_18_V_read_8_reg_9874_pp0_iter4_reg;
        data_18_V_read_8_reg_9874_pp0_iter6_reg <= data_18_V_read_8_reg_9874_pp0_iter5_reg;
        data_19_V_read_8_reg_9845 <= data_19_V_read_int_reg;
        data_19_V_read_8_reg_9845_pp0_iter1_reg <= data_19_V_read_8_reg_9845;
        data_19_V_read_8_reg_9845_pp0_iter2_reg <= data_19_V_read_8_reg_9845_pp0_iter1_reg;
        data_19_V_read_8_reg_9845_pp0_iter3_reg <= data_19_V_read_8_reg_9845_pp0_iter2_reg;
        data_19_V_read_8_reg_9845_pp0_iter4_reg <= data_19_V_read_8_reg_9845_pp0_iter3_reg;
        data_19_V_read_8_reg_9845_pp0_iter5_reg <= data_19_V_read_8_reg_9845_pp0_iter4_reg;
        data_19_V_read_8_reg_9845_pp0_iter6_reg <= data_19_V_read_8_reg_9845_pp0_iter5_reg;
        data_1_V_read_10_reg_10323 <= data_1_V_read_int_reg;
        data_20_V_read21_reg_9814 <= data_20_V_read_int_reg;
        data_20_V_read21_reg_9814_pp0_iter1_reg <= data_20_V_read21_reg_9814;
        data_20_V_read21_reg_9814_pp0_iter2_reg <= data_20_V_read21_reg_9814_pp0_iter1_reg;
        data_20_V_read21_reg_9814_pp0_iter3_reg <= data_20_V_read21_reg_9814_pp0_iter2_reg;
        data_20_V_read21_reg_9814_pp0_iter4_reg <= data_20_V_read21_reg_9814_pp0_iter3_reg;
        data_20_V_read21_reg_9814_pp0_iter5_reg <= data_20_V_read21_reg_9814_pp0_iter4_reg;
        data_20_V_read21_reg_9814_pp0_iter6_reg <= data_20_V_read21_reg_9814_pp0_iter5_reg;
        data_20_V_read21_reg_9814_pp0_iter7_reg <= data_20_V_read21_reg_9814_pp0_iter6_reg;
        data_21_V_read22_reg_9784 <= data_21_V_read_int_reg;
        data_21_V_read22_reg_9784_pp0_iter1_reg <= data_21_V_read22_reg_9784;
        data_21_V_read22_reg_9784_pp0_iter2_reg <= data_21_V_read22_reg_9784_pp0_iter1_reg;
        data_21_V_read22_reg_9784_pp0_iter3_reg <= data_21_V_read22_reg_9784_pp0_iter2_reg;
        data_21_V_read22_reg_9784_pp0_iter4_reg <= data_21_V_read22_reg_9784_pp0_iter3_reg;
        data_21_V_read22_reg_9784_pp0_iter5_reg <= data_21_V_read22_reg_9784_pp0_iter4_reg;
        data_21_V_read22_reg_9784_pp0_iter6_reg <= data_21_V_read22_reg_9784_pp0_iter5_reg;
        data_21_V_read22_reg_9784_pp0_iter7_reg <= data_21_V_read22_reg_9784_pp0_iter6_reg;
        data_22_V_read23_reg_9756 <= data_22_V_read_int_reg;
        data_22_V_read23_reg_9756_pp0_iter1_reg <= data_22_V_read23_reg_9756;
        data_22_V_read23_reg_9756_pp0_iter2_reg <= data_22_V_read23_reg_9756_pp0_iter1_reg;
        data_22_V_read23_reg_9756_pp0_iter3_reg <= data_22_V_read23_reg_9756_pp0_iter2_reg;
        data_22_V_read23_reg_9756_pp0_iter4_reg <= data_22_V_read23_reg_9756_pp0_iter3_reg;
        data_22_V_read23_reg_9756_pp0_iter5_reg <= data_22_V_read23_reg_9756_pp0_iter4_reg;
        data_22_V_read23_reg_9756_pp0_iter6_reg <= data_22_V_read23_reg_9756_pp0_iter5_reg;
        data_22_V_read23_reg_9756_pp0_iter7_reg <= data_22_V_read23_reg_9756_pp0_iter6_reg;
        data_22_V_read23_reg_9756_pp0_iter8_reg <= data_22_V_read23_reg_9756_pp0_iter7_reg;
        data_23_V_read24_reg_9730 <= data_23_V_read_int_reg;
        data_23_V_read24_reg_9730_pp0_iter1_reg <= data_23_V_read24_reg_9730;
        data_23_V_read24_reg_9730_pp0_iter2_reg <= data_23_V_read24_reg_9730_pp0_iter1_reg;
        data_23_V_read24_reg_9730_pp0_iter3_reg <= data_23_V_read24_reg_9730_pp0_iter2_reg;
        data_23_V_read24_reg_9730_pp0_iter4_reg <= data_23_V_read24_reg_9730_pp0_iter3_reg;
        data_23_V_read24_reg_9730_pp0_iter5_reg <= data_23_V_read24_reg_9730_pp0_iter4_reg;
        data_23_V_read24_reg_9730_pp0_iter6_reg <= data_23_V_read24_reg_9730_pp0_iter5_reg;
        data_23_V_read24_reg_9730_pp0_iter7_reg <= data_23_V_read24_reg_9730_pp0_iter6_reg;
        data_24_V_read25_reg_9704 <= data_24_V_read_int_reg;
        data_24_V_read25_reg_9704_pp0_iter1_reg <= data_24_V_read25_reg_9704;
        data_24_V_read25_reg_9704_pp0_iter2_reg <= data_24_V_read25_reg_9704_pp0_iter1_reg;
        data_24_V_read25_reg_9704_pp0_iter3_reg <= data_24_V_read25_reg_9704_pp0_iter2_reg;
        data_24_V_read25_reg_9704_pp0_iter4_reg <= data_24_V_read25_reg_9704_pp0_iter3_reg;
        data_24_V_read25_reg_9704_pp0_iter5_reg <= data_24_V_read25_reg_9704_pp0_iter4_reg;
        data_24_V_read25_reg_9704_pp0_iter6_reg <= data_24_V_read25_reg_9704_pp0_iter5_reg;
        data_24_V_read25_reg_9704_pp0_iter7_reg <= data_24_V_read25_reg_9704_pp0_iter6_reg;
        data_24_V_read25_reg_9704_pp0_iter8_reg <= data_24_V_read25_reg_9704_pp0_iter7_reg;
        data_25_V_read26_reg_9677 <= data_25_V_read_int_reg;
        data_25_V_read26_reg_9677_pp0_iter1_reg <= data_25_V_read26_reg_9677;
        data_25_V_read26_reg_9677_pp0_iter2_reg <= data_25_V_read26_reg_9677_pp0_iter1_reg;
        data_25_V_read26_reg_9677_pp0_iter3_reg <= data_25_V_read26_reg_9677_pp0_iter2_reg;
        data_25_V_read26_reg_9677_pp0_iter4_reg <= data_25_V_read26_reg_9677_pp0_iter3_reg;
        data_25_V_read26_reg_9677_pp0_iter5_reg <= data_25_V_read26_reg_9677_pp0_iter4_reg;
        data_25_V_read26_reg_9677_pp0_iter6_reg <= data_25_V_read26_reg_9677_pp0_iter5_reg;
        data_25_V_read26_reg_9677_pp0_iter7_reg <= data_25_V_read26_reg_9677_pp0_iter6_reg;
        data_25_V_read26_reg_9677_pp0_iter8_reg <= data_25_V_read26_reg_9677_pp0_iter7_reg;
        data_26_V_read27_reg_9652 <= data_26_V_read_int_reg;
        data_26_V_read27_reg_9652_pp0_iter1_reg <= data_26_V_read27_reg_9652;
        data_26_V_read27_reg_9652_pp0_iter2_reg <= data_26_V_read27_reg_9652_pp0_iter1_reg;
        data_26_V_read27_reg_9652_pp0_iter3_reg <= data_26_V_read27_reg_9652_pp0_iter2_reg;
        data_26_V_read27_reg_9652_pp0_iter4_reg <= data_26_V_read27_reg_9652_pp0_iter3_reg;
        data_26_V_read27_reg_9652_pp0_iter5_reg <= data_26_V_read27_reg_9652_pp0_iter4_reg;
        data_26_V_read27_reg_9652_pp0_iter6_reg <= data_26_V_read27_reg_9652_pp0_iter5_reg;
        data_26_V_read27_reg_9652_pp0_iter7_reg <= data_26_V_read27_reg_9652_pp0_iter6_reg;
        data_26_V_read27_reg_9652_pp0_iter8_reg <= data_26_V_read27_reg_9652_pp0_iter7_reg;
        data_27_V_read28_reg_9625 <= data_27_V_read_int_reg;
        data_27_V_read28_reg_9625_pp0_iter1_reg <= data_27_V_read28_reg_9625;
        data_27_V_read28_reg_9625_pp0_iter2_reg <= data_27_V_read28_reg_9625_pp0_iter1_reg;
        data_27_V_read28_reg_9625_pp0_iter3_reg <= data_27_V_read28_reg_9625_pp0_iter2_reg;
        data_27_V_read28_reg_9625_pp0_iter4_reg <= data_27_V_read28_reg_9625_pp0_iter3_reg;
        data_27_V_read28_reg_9625_pp0_iter5_reg <= data_27_V_read28_reg_9625_pp0_iter4_reg;
        data_27_V_read28_reg_9625_pp0_iter6_reg <= data_27_V_read28_reg_9625_pp0_iter5_reg;
        data_27_V_read28_reg_9625_pp0_iter7_reg <= data_27_V_read28_reg_9625_pp0_iter6_reg;
        data_27_V_read28_reg_9625_pp0_iter8_reg <= data_27_V_read28_reg_9625_pp0_iter7_reg;
        data_28_V_read_8_reg_9598 <= data_28_V_read_int_reg;
        data_28_V_read_8_reg_9598_pp0_iter1_reg <= data_28_V_read_8_reg_9598;
        data_28_V_read_8_reg_9598_pp0_iter2_reg <= data_28_V_read_8_reg_9598_pp0_iter1_reg;
        data_28_V_read_8_reg_9598_pp0_iter3_reg <= data_28_V_read_8_reg_9598_pp0_iter2_reg;
        data_28_V_read_8_reg_9598_pp0_iter4_reg <= data_28_V_read_8_reg_9598_pp0_iter3_reg;
        data_28_V_read_8_reg_9598_pp0_iter5_reg <= data_28_V_read_8_reg_9598_pp0_iter4_reg;
        data_28_V_read_8_reg_9598_pp0_iter6_reg <= data_28_V_read_8_reg_9598_pp0_iter5_reg;
        data_28_V_read_8_reg_9598_pp0_iter7_reg <= data_28_V_read_8_reg_9598_pp0_iter6_reg;
        data_28_V_read_8_reg_9598_pp0_iter8_reg <= data_28_V_read_8_reg_9598_pp0_iter7_reg;
        data_29_V_read_8_reg_9573 <= data_29_V_read_int_reg;
        data_29_V_read_8_reg_9573_pp0_iter1_reg <= data_29_V_read_8_reg_9573;
        data_29_V_read_8_reg_9573_pp0_iter2_reg <= data_29_V_read_8_reg_9573_pp0_iter1_reg;
        data_29_V_read_8_reg_9573_pp0_iter3_reg <= data_29_V_read_8_reg_9573_pp0_iter2_reg;
        data_29_V_read_8_reg_9573_pp0_iter4_reg <= data_29_V_read_8_reg_9573_pp0_iter3_reg;
        data_29_V_read_8_reg_9573_pp0_iter5_reg <= data_29_V_read_8_reg_9573_pp0_iter4_reg;
        data_29_V_read_8_reg_9573_pp0_iter6_reg <= data_29_V_read_8_reg_9573_pp0_iter5_reg;
        data_29_V_read_8_reg_9573_pp0_iter7_reg <= data_29_V_read_8_reg_9573_pp0_iter6_reg;
        data_29_V_read_8_reg_9573_pp0_iter8_reg <= data_29_V_read_8_reg_9573_pp0_iter7_reg;
        data_29_V_read_8_reg_9573_pp0_iter9_reg <= data_29_V_read_8_reg_9573_pp0_iter8_reg;
        data_2_V_read_10_reg_10312 <= data_2_V_read_int_reg;
        data_2_V_read_10_reg_10312_pp0_iter1_reg <= data_2_V_read_10_reg_10312;
        data_30_V_read31_reg_9549 <= data_30_V_read_int_reg;
        data_30_V_read31_reg_9549_pp0_iter1_reg <= data_30_V_read31_reg_9549;
        data_30_V_read31_reg_9549_pp0_iter2_reg <= data_30_V_read31_reg_9549_pp0_iter1_reg;
        data_30_V_read31_reg_9549_pp0_iter3_reg <= data_30_V_read31_reg_9549_pp0_iter2_reg;
        data_30_V_read31_reg_9549_pp0_iter4_reg <= data_30_V_read31_reg_9549_pp0_iter3_reg;
        data_30_V_read31_reg_9549_pp0_iter5_reg <= data_30_V_read31_reg_9549_pp0_iter4_reg;
        data_30_V_read31_reg_9549_pp0_iter6_reg <= data_30_V_read31_reg_9549_pp0_iter5_reg;
        data_30_V_read31_reg_9549_pp0_iter7_reg <= data_30_V_read31_reg_9549_pp0_iter6_reg;
        data_30_V_read31_reg_9549_pp0_iter8_reg <= data_30_V_read31_reg_9549_pp0_iter7_reg;
        data_30_V_read31_reg_9549_pp0_iter9_reg <= data_30_V_read31_reg_9549_pp0_iter8_reg;
        data_31_V_read32_reg_9521 <= data_31_V_read_int_reg;
        data_31_V_read32_reg_9521_pp0_iter1_reg <= data_31_V_read32_reg_9521;
        data_31_V_read32_reg_9521_pp0_iter2_reg <= data_31_V_read32_reg_9521_pp0_iter1_reg;
        data_31_V_read32_reg_9521_pp0_iter3_reg <= data_31_V_read32_reg_9521_pp0_iter2_reg;
        data_31_V_read32_reg_9521_pp0_iter4_reg <= data_31_V_read32_reg_9521_pp0_iter3_reg;
        data_31_V_read32_reg_9521_pp0_iter5_reg <= data_31_V_read32_reg_9521_pp0_iter4_reg;
        data_31_V_read32_reg_9521_pp0_iter6_reg <= data_31_V_read32_reg_9521_pp0_iter5_reg;
        data_31_V_read32_reg_9521_pp0_iter7_reg <= data_31_V_read32_reg_9521_pp0_iter6_reg;
        data_31_V_read32_reg_9521_pp0_iter8_reg <= data_31_V_read32_reg_9521_pp0_iter7_reg;
        data_31_V_read32_reg_9521_pp0_iter9_reg <= data_31_V_read32_reg_9521_pp0_iter8_reg;
        data_32_V_read_3_reg_9492 <= data_32_V_read_int_reg;
        data_32_V_read_3_reg_9492_pp0_iter1_reg <= data_32_V_read_3_reg_9492;
        data_32_V_read_3_reg_9492_pp0_iter2_reg <= data_32_V_read_3_reg_9492_pp0_iter1_reg;
        data_32_V_read_3_reg_9492_pp0_iter3_reg <= data_32_V_read_3_reg_9492_pp0_iter2_reg;
        data_32_V_read_3_reg_9492_pp0_iter4_reg <= data_32_V_read_3_reg_9492_pp0_iter3_reg;
        data_32_V_read_3_reg_9492_pp0_iter5_reg <= data_32_V_read_3_reg_9492_pp0_iter4_reg;
        data_32_V_read_3_reg_9492_pp0_iter6_reg <= data_32_V_read_3_reg_9492_pp0_iter5_reg;
        data_32_V_read_3_reg_9492_pp0_iter7_reg <= data_32_V_read_3_reg_9492_pp0_iter6_reg;
        data_32_V_read_3_reg_9492_pp0_iter8_reg <= data_32_V_read_3_reg_9492_pp0_iter7_reg;
        data_32_V_read_3_reg_9492_pp0_iter9_reg <= data_32_V_read_3_reg_9492_pp0_iter8_reg;
        data_33_V_read_3_reg_9463 <= data_33_V_read_int_reg;
        data_33_V_read_3_reg_9463_pp0_iter10_reg <= data_33_V_read_3_reg_9463_pp0_iter9_reg;
        data_33_V_read_3_reg_9463_pp0_iter1_reg <= data_33_V_read_3_reg_9463;
        data_33_V_read_3_reg_9463_pp0_iter2_reg <= data_33_V_read_3_reg_9463_pp0_iter1_reg;
        data_33_V_read_3_reg_9463_pp0_iter3_reg <= data_33_V_read_3_reg_9463_pp0_iter2_reg;
        data_33_V_read_3_reg_9463_pp0_iter4_reg <= data_33_V_read_3_reg_9463_pp0_iter3_reg;
        data_33_V_read_3_reg_9463_pp0_iter5_reg <= data_33_V_read_3_reg_9463_pp0_iter4_reg;
        data_33_V_read_3_reg_9463_pp0_iter6_reg <= data_33_V_read_3_reg_9463_pp0_iter5_reg;
        data_33_V_read_3_reg_9463_pp0_iter7_reg <= data_33_V_read_3_reg_9463_pp0_iter6_reg;
        data_33_V_read_3_reg_9463_pp0_iter8_reg <= data_33_V_read_3_reg_9463_pp0_iter7_reg;
        data_33_V_read_3_reg_9463_pp0_iter9_reg <= data_33_V_read_3_reg_9463_pp0_iter8_reg;
        data_34_V_read_3_reg_9434 <= data_34_V_read_int_reg;
        data_34_V_read_3_reg_9434_pp0_iter10_reg <= data_34_V_read_3_reg_9434_pp0_iter9_reg;
        data_34_V_read_3_reg_9434_pp0_iter1_reg <= data_34_V_read_3_reg_9434;
        data_34_V_read_3_reg_9434_pp0_iter2_reg <= data_34_V_read_3_reg_9434_pp0_iter1_reg;
        data_34_V_read_3_reg_9434_pp0_iter3_reg <= data_34_V_read_3_reg_9434_pp0_iter2_reg;
        data_34_V_read_3_reg_9434_pp0_iter4_reg <= data_34_V_read_3_reg_9434_pp0_iter3_reg;
        data_34_V_read_3_reg_9434_pp0_iter5_reg <= data_34_V_read_3_reg_9434_pp0_iter4_reg;
        data_34_V_read_3_reg_9434_pp0_iter6_reg <= data_34_V_read_3_reg_9434_pp0_iter5_reg;
        data_34_V_read_3_reg_9434_pp0_iter7_reg <= data_34_V_read_3_reg_9434_pp0_iter6_reg;
        data_34_V_read_3_reg_9434_pp0_iter8_reg <= data_34_V_read_3_reg_9434_pp0_iter7_reg;
        data_34_V_read_3_reg_9434_pp0_iter9_reg <= data_34_V_read_3_reg_9434_pp0_iter8_reg;
        data_35_V_read_3_reg_9410 <= data_35_V_read_int_reg;
        data_35_V_read_3_reg_9410_pp0_iter10_reg <= data_35_V_read_3_reg_9410_pp0_iter9_reg;
        data_35_V_read_3_reg_9410_pp0_iter1_reg <= data_35_V_read_3_reg_9410;
        data_35_V_read_3_reg_9410_pp0_iter2_reg <= data_35_V_read_3_reg_9410_pp0_iter1_reg;
        data_35_V_read_3_reg_9410_pp0_iter3_reg <= data_35_V_read_3_reg_9410_pp0_iter2_reg;
        data_35_V_read_3_reg_9410_pp0_iter4_reg <= data_35_V_read_3_reg_9410_pp0_iter3_reg;
        data_35_V_read_3_reg_9410_pp0_iter5_reg <= data_35_V_read_3_reg_9410_pp0_iter4_reg;
        data_35_V_read_3_reg_9410_pp0_iter6_reg <= data_35_V_read_3_reg_9410_pp0_iter5_reg;
        data_35_V_read_3_reg_9410_pp0_iter7_reg <= data_35_V_read_3_reg_9410_pp0_iter6_reg;
        data_35_V_read_3_reg_9410_pp0_iter8_reg <= data_35_V_read_3_reg_9410_pp0_iter7_reg;
        data_35_V_read_3_reg_9410_pp0_iter9_reg <= data_35_V_read_3_reg_9410_pp0_iter8_reg;
        data_36_V_read_3_reg_9383 <= data_36_V_read_int_reg;
        data_36_V_read_3_reg_9383_pp0_iter10_reg <= data_36_V_read_3_reg_9383_pp0_iter9_reg;
        data_36_V_read_3_reg_9383_pp0_iter1_reg <= data_36_V_read_3_reg_9383;
        data_36_V_read_3_reg_9383_pp0_iter2_reg <= data_36_V_read_3_reg_9383_pp0_iter1_reg;
        data_36_V_read_3_reg_9383_pp0_iter3_reg <= data_36_V_read_3_reg_9383_pp0_iter2_reg;
        data_36_V_read_3_reg_9383_pp0_iter4_reg <= data_36_V_read_3_reg_9383_pp0_iter3_reg;
        data_36_V_read_3_reg_9383_pp0_iter5_reg <= data_36_V_read_3_reg_9383_pp0_iter4_reg;
        data_36_V_read_3_reg_9383_pp0_iter6_reg <= data_36_V_read_3_reg_9383_pp0_iter5_reg;
        data_36_V_read_3_reg_9383_pp0_iter7_reg <= data_36_V_read_3_reg_9383_pp0_iter6_reg;
        data_36_V_read_3_reg_9383_pp0_iter8_reg <= data_36_V_read_3_reg_9383_pp0_iter7_reg;
        data_36_V_read_3_reg_9383_pp0_iter9_reg <= data_36_V_read_3_reg_9383_pp0_iter8_reg;
        data_37_V_read_3_reg_9353 <= data_37_V_read_int_reg;
        data_37_V_read_3_reg_9353_pp0_iter10_reg <= data_37_V_read_3_reg_9353_pp0_iter9_reg;
        data_37_V_read_3_reg_9353_pp0_iter1_reg <= data_37_V_read_3_reg_9353;
        data_37_V_read_3_reg_9353_pp0_iter2_reg <= data_37_V_read_3_reg_9353_pp0_iter1_reg;
        data_37_V_read_3_reg_9353_pp0_iter3_reg <= data_37_V_read_3_reg_9353_pp0_iter2_reg;
        data_37_V_read_3_reg_9353_pp0_iter4_reg <= data_37_V_read_3_reg_9353_pp0_iter3_reg;
        data_37_V_read_3_reg_9353_pp0_iter5_reg <= data_37_V_read_3_reg_9353_pp0_iter4_reg;
        data_37_V_read_3_reg_9353_pp0_iter6_reg <= data_37_V_read_3_reg_9353_pp0_iter5_reg;
        data_37_V_read_3_reg_9353_pp0_iter7_reg <= data_37_V_read_3_reg_9353_pp0_iter6_reg;
        data_37_V_read_3_reg_9353_pp0_iter8_reg <= data_37_V_read_3_reg_9353_pp0_iter7_reg;
        data_37_V_read_3_reg_9353_pp0_iter9_reg <= data_37_V_read_3_reg_9353_pp0_iter8_reg;
        data_38_V_read_3_reg_9328 <= data_38_V_read_int_reg;
        data_38_V_read_3_reg_9328_pp0_iter10_reg <= data_38_V_read_3_reg_9328_pp0_iter9_reg;
        data_38_V_read_3_reg_9328_pp0_iter11_reg <= data_38_V_read_3_reg_9328_pp0_iter10_reg;
        data_38_V_read_3_reg_9328_pp0_iter1_reg <= data_38_V_read_3_reg_9328;
        data_38_V_read_3_reg_9328_pp0_iter2_reg <= data_38_V_read_3_reg_9328_pp0_iter1_reg;
        data_38_V_read_3_reg_9328_pp0_iter3_reg <= data_38_V_read_3_reg_9328_pp0_iter2_reg;
        data_38_V_read_3_reg_9328_pp0_iter4_reg <= data_38_V_read_3_reg_9328_pp0_iter3_reg;
        data_38_V_read_3_reg_9328_pp0_iter5_reg <= data_38_V_read_3_reg_9328_pp0_iter4_reg;
        data_38_V_read_3_reg_9328_pp0_iter6_reg <= data_38_V_read_3_reg_9328_pp0_iter5_reg;
        data_38_V_read_3_reg_9328_pp0_iter7_reg <= data_38_V_read_3_reg_9328_pp0_iter6_reg;
        data_38_V_read_3_reg_9328_pp0_iter8_reg <= data_38_V_read_3_reg_9328_pp0_iter7_reg;
        data_38_V_read_3_reg_9328_pp0_iter9_reg <= data_38_V_read_3_reg_9328_pp0_iter8_reg;
        data_39_V_read_3_reg_9301 <= data_39_V_read_int_reg;
        data_39_V_read_3_reg_9301_pp0_iter10_reg <= data_39_V_read_3_reg_9301_pp0_iter9_reg;
        data_39_V_read_3_reg_9301_pp0_iter11_reg <= data_39_V_read_3_reg_9301_pp0_iter10_reg;
        data_39_V_read_3_reg_9301_pp0_iter1_reg <= data_39_V_read_3_reg_9301;
        data_39_V_read_3_reg_9301_pp0_iter2_reg <= data_39_V_read_3_reg_9301_pp0_iter1_reg;
        data_39_V_read_3_reg_9301_pp0_iter3_reg <= data_39_V_read_3_reg_9301_pp0_iter2_reg;
        data_39_V_read_3_reg_9301_pp0_iter4_reg <= data_39_V_read_3_reg_9301_pp0_iter3_reg;
        data_39_V_read_3_reg_9301_pp0_iter5_reg <= data_39_V_read_3_reg_9301_pp0_iter4_reg;
        data_39_V_read_3_reg_9301_pp0_iter6_reg <= data_39_V_read_3_reg_9301_pp0_iter5_reg;
        data_39_V_read_3_reg_9301_pp0_iter7_reg <= data_39_V_read_3_reg_9301_pp0_iter6_reg;
        data_39_V_read_3_reg_9301_pp0_iter8_reg <= data_39_V_read_3_reg_9301_pp0_iter7_reg;
        data_39_V_read_3_reg_9301_pp0_iter9_reg <= data_39_V_read_3_reg_9301_pp0_iter8_reg;
        data_3_V_read_10_reg_10295 <= data_3_V_read_int_reg;
        data_3_V_read_10_reg_10295_pp0_iter1_reg <= data_3_V_read_10_reg_10295;
        data_3_V_read_10_reg_10295_pp0_iter2_reg <= data_3_V_read_10_reg_10295_pp0_iter1_reg;
        data_40_V_read41_reg_9272 <= data_40_V_read_int_reg;
        data_40_V_read41_reg_9272_pp0_iter10_reg <= data_40_V_read41_reg_9272_pp0_iter9_reg;
        data_40_V_read41_reg_9272_pp0_iter11_reg <= data_40_V_read41_reg_9272_pp0_iter10_reg;
        data_40_V_read41_reg_9272_pp0_iter1_reg <= data_40_V_read41_reg_9272;
        data_40_V_read41_reg_9272_pp0_iter2_reg <= data_40_V_read41_reg_9272_pp0_iter1_reg;
        data_40_V_read41_reg_9272_pp0_iter3_reg <= data_40_V_read41_reg_9272_pp0_iter2_reg;
        data_40_V_read41_reg_9272_pp0_iter4_reg <= data_40_V_read41_reg_9272_pp0_iter3_reg;
        data_40_V_read41_reg_9272_pp0_iter5_reg <= data_40_V_read41_reg_9272_pp0_iter4_reg;
        data_40_V_read41_reg_9272_pp0_iter6_reg <= data_40_V_read41_reg_9272_pp0_iter5_reg;
        data_40_V_read41_reg_9272_pp0_iter7_reg <= data_40_V_read41_reg_9272_pp0_iter6_reg;
        data_40_V_read41_reg_9272_pp0_iter8_reg <= data_40_V_read41_reg_9272_pp0_iter7_reg;
        data_40_V_read41_reg_9272_pp0_iter9_reg <= data_40_V_read41_reg_9272_pp0_iter8_reg;
        data_41_V_read42_reg_9242 <= data_41_V_read_int_reg;
        data_41_V_read42_reg_9242_pp0_iter10_reg <= data_41_V_read42_reg_9242_pp0_iter9_reg;
        data_41_V_read42_reg_9242_pp0_iter11_reg <= data_41_V_read42_reg_9242_pp0_iter10_reg;
        data_41_V_read42_reg_9242_pp0_iter1_reg <= data_41_V_read42_reg_9242;
        data_41_V_read42_reg_9242_pp0_iter2_reg <= data_41_V_read42_reg_9242_pp0_iter1_reg;
        data_41_V_read42_reg_9242_pp0_iter3_reg <= data_41_V_read42_reg_9242_pp0_iter2_reg;
        data_41_V_read42_reg_9242_pp0_iter4_reg <= data_41_V_read42_reg_9242_pp0_iter3_reg;
        data_41_V_read42_reg_9242_pp0_iter5_reg <= data_41_V_read42_reg_9242_pp0_iter4_reg;
        data_41_V_read42_reg_9242_pp0_iter6_reg <= data_41_V_read42_reg_9242_pp0_iter5_reg;
        data_41_V_read42_reg_9242_pp0_iter7_reg <= data_41_V_read42_reg_9242_pp0_iter6_reg;
        data_41_V_read42_reg_9242_pp0_iter8_reg <= data_41_V_read42_reg_9242_pp0_iter7_reg;
        data_41_V_read42_reg_9242_pp0_iter9_reg <= data_41_V_read42_reg_9242_pp0_iter8_reg;
        data_42_V_read_3_reg_9212 <= data_42_V_read_int_reg;
        data_42_V_read_3_reg_9212_pp0_iter10_reg <= data_42_V_read_3_reg_9212_pp0_iter9_reg;
        data_42_V_read_3_reg_9212_pp0_iter11_reg <= data_42_V_read_3_reg_9212_pp0_iter10_reg;
        data_42_V_read_3_reg_9212_pp0_iter12_reg <= data_42_V_read_3_reg_9212_pp0_iter11_reg;
        data_42_V_read_3_reg_9212_pp0_iter1_reg <= data_42_V_read_3_reg_9212;
        data_42_V_read_3_reg_9212_pp0_iter2_reg <= data_42_V_read_3_reg_9212_pp0_iter1_reg;
        data_42_V_read_3_reg_9212_pp0_iter3_reg <= data_42_V_read_3_reg_9212_pp0_iter2_reg;
        data_42_V_read_3_reg_9212_pp0_iter4_reg <= data_42_V_read_3_reg_9212_pp0_iter3_reg;
        data_42_V_read_3_reg_9212_pp0_iter5_reg <= data_42_V_read_3_reg_9212_pp0_iter4_reg;
        data_42_V_read_3_reg_9212_pp0_iter6_reg <= data_42_V_read_3_reg_9212_pp0_iter5_reg;
        data_42_V_read_3_reg_9212_pp0_iter7_reg <= data_42_V_read_3_reg_9212_pp0_iter6_reg;
        data_42_V_read_3_reg_9212_pp0_iter8_reg <= data_42_V_read_3_reg_9212_pp0_iter7_reg;
        data_42_V_read_3_reg_9212_pp0_iter9_reg <= data_42_V_read_3_reg_9212_pp0_iter8_reg;
        data_43_V_read_3_reg_9184 <= data_43_V_read_int_reg;
        data_43_V_read_3_reg_9184_pp0_iter10_reg <= data_43_V_read_3_reg_9184_pp0_iter9_reg;
        data_43_V_read_3_reg_9184_pp0_iter11_reg <= data_43_V_read_3_reg_9184_pp0_iter10_reg;
        data_43_V_read_3_reg_9184_pp0_iter12_reg <= data_43_V_read_3_reg_9184_pp0_iter11_reg;
        data_43_V_read_3_reg_9184_pp0_iter1_reg <= data_43_V_read_3_reg_9184;
        data_43_V_read_3_reg_9184_pp0_iter2_reg <= data_43_V_read_3_reg_9184_pp0_iter1_reg;
        data_43_V_read_3_reg_9184_pp0_iter3_reg <= data_43_V_read_3_reg_9184_pp0_iter2_reg;
        data_43_V_read_3_reg_9184_pp0_iter4_reg <= data_43_V_read_3_reg_9184_pp0_iter3_reg;
        data_43_V_read_3_reg_9184_pp0_iter5_reg <= data_43_V_read_3_reg_9184_pp0_iter4_reg;
        data_43_V_read_3_reg_9184_pp0_iter6_reg <= data_43_V_read_3_reg_9184_pp0_iter5_reg;
        data_43_V_read_3_reg_9184_pp0_iter7_reg <= data_43_V_read_3_reg_9184_pp0_iter6_reg;
        data_43_V_read_3_reg_9184_pp0_iter8_reg <= data_43_V_read_3_reg_9184_pp0_iter7_reg;
        data_43_V_read_3_reg_9184_pp0_iter9_reg <= data_43_V_read_3_reg_9184_pp0_iter8_reg;
        data_44_V_read_3_reg_9154 <= data_44_V_read_int_reg;
        data_44_V_read_3_reg_9154_pp0_iter10_reg <= data_44_V_read_3_reg_9154_pp0_iter9_reg;
        data_44_V_read_3_reg_9154_pp0_iter11_reg <= data_44_V_read_3_reg_9154_pp0_iter10_reg;
        data_44_V_read_3_reg_9154_pp0_iter12_reg <= data_44_V_read_3_reg_9154_pp0_iter11_reg;
        data_44_V_read_3_reg_9154_pp0_iter1_reg <= data_44_V_read_3_reg_9154;
        data_44_V_read_3_reg_9154_pp0_iter2_reg <= data_44_V_read_3_reg_9154_pp0_iter1_reg;
        data_44_V_read_3_reg_9154_pp0_iter3_reg <= data_44_V_read_3_reg_9154_pp0_iter2_reg;
        data_44_V_read_3_reg_9154_pp0_iter4_reg <= data_44_V_read_3_reg_9154_pp0_iter3_reg;
        data_44_V_read_3_reg_9154_pp0_iter5_reg <= data_44_V_read_3_reg_9154_pp0_iter4_reg;
        data_44_V_read_3_reg_9154_pp0_iter6_reg <= data_44_V_read_3_reg_9154_pp0_iter5_reg;
        data_44_V_read_3_reg_9154_pp0_iter7_reg <= data_44_V_read_3_reg_9154_pp0_iter6_reg;
        data_44_V_read_3_reg_9154_pp0_iter8_reg <= data_44_V_read_3_reg_9154_pp0_iter7_reg;
        data_44_V_read_3_reg_9154_pp0_iter9_reg <= data_44_V_read_3_reg_9154_pp0_iter8_reg;
        data_45_V_read_3_reg_9125 <= data_45_V_read_int_reg;
        data_45_V_read_3_reg_9125_pp0_iter10_reg <= data_45_V_read_3_reg_9125_pp0_iter9_reg;
        data_45_V_read_3_reg_9125_pp0_iter11_reg <= data_45_V_read_3_reg_9125_pp0_iter10_reg;
        data_45_V_read_3_reg_9125_pp0_iter12_reg <= data_45_V_read_3_reg_9125_pp0_iter11_reg;
        data_45_V_read_3_reg_9125_pp0_iter1_reg <= data_45_V_read_3_reg_9125;
        data_45_V_read_3_reg_9125_pp0_iter2_reg <= data_45_V_read_3_reg_9125_pp0_iter1_reg;
        data_45_V_read_3_reg_9125_pp0_iter3_reg <= data_45_V_read_3_reg_9125_pp0_iter2_reg;
        data_45_V_read_3_reg_9125_pp0_iter4_reg <= data_45_V_read_3_reg_9125_pp0_iter3_reg;
        data_45_V_read_3_reg_9125_pp0_iter5_reg <= data_45_V_read_3_reg_9125_pp0_iter4_reg;
        data_45_V_read_3_reg_9125_pp0_iter6_reg <= data_45_V_read_3_reg_9125_pp0_iter5_reg;
        data_45_V_read_3_reg_9125_pp0_iter7_reg <= data_45_V_read_3_reg_9125_pp0_iter6_reg;
        data_45_V_read_3_reg_9125_pp0_iter8_reg <= data_45_V_read_3_reg_9125_pp0_iter7_reg;
        data_45_V_read_3_reg_9125_pp0_iter9_reg <= data_45_V_read_3_reg_9125_pp0_iter8_reg;
        data_46_V_read_3_reg_9094 <= data_46_V_read_int_reg;
        data_46_V_read_3_reg_9094_pp0_iter10_reg <= data_46_V_read_3_reg_9094_pp0_iter9_reg;
        data_46_V_read_3_reg_9094_pp0_iter11_reg <= data_46_V_read_3_reg_9094_pp0_iter10_reg;
        data_46_V_read_3_reg_9094_pp0_iter12_reg <= data_46_V_read_3_reg_9094_pp0_iter11_reg;
        data_46_V_read_3_reg_9094_pp0_iter13_reg <= data_46_V_read_3_reg_9094_pp0_iter12_reg;
        data_46_V_read_3_reg_9094_pp0_iter1_reg <= data_46_V_read_3_reg_9094;
        data_46_V_read_3_reg_9094_pp0_iter2_reg <= data_46_V_read_3_reg_9094_pp0_iter1_reg;
        data_46_V_read_3_reg_9094_pp0_iter3_reg <= data_46_V_read_3_reg_9094_pp0_iter2_reg;
        data_46_V_read_3_reg_9094_pp0_iter4_reg <= data_46_V_read_3_reg_9094_pp0_iter3_reg;
        data_46_V_read_3_reg_9094_pp0_iter5_reg <= data_46_V_read_3_reg_9094_pp0_iter4_reg;
        data_46_V_read_3_reg_9094_pp0_iter6_reg <= data_46_V_read_3_reg_9094_pp0_iter5_reg;
        data_46_V_read_3_reg_9094_pp0_iter7_reg <= data_46_V_read_3_reg_9094_pp0_iter6_reg;
        data_46_V_read_3_reg_9094_pp0_iter8_reg <= data_46_V_read_3_reg_9094_pp0_iter7_reg;
        data_46_V_read_3_reg_9094_pp0_iter9_reg <= data_46_V_read_3_reg_9094_pp0_iter8_reg;
        data_47_V_read_3_reg_9066 <= data_47_V_read_int_reg;
        data_47_V_read_3_reg_9066_pp0_iter10_reg <= data_47_V_read_3_reg_9066_pp0_iter9_reg;
        data_47_V_read_3_reg_9066_pp0_iter11_reg <= data_47_V_read_3_reg_9066_pp0_iter10_reg;
        data_47_V_read_3_reg_9066_pp0_iter12_reg <= data_47_V_read_3_reg_9066_pp0_iter11_reg;
        data_47_V_read_3_reg_9066_pp0_iter13_reg <= data_47_V_read_3_reg_9066_pp0_iter12_reg;
        data_47_V_read_3_reg_9066_pp0_iter1_reg <= data_47_V_read_3_reg_9066;
        data_47_V_read_3_reg_9066_pp0_iter2_reg <= data_47_V_read_3_reg_9066_pp0_iter1_reg;
        data_47_V_read_3_reg_9066_pp0_iter3_reg <= data_47_V_read_3_reg_9066_pp0_iter2_reg;
        data_47_V_read_3_reg_9066_pp0_iter4_reg <= data_47_V_read_3_reg_9066_pp0_iter3_reg;
        data_47_V_read_3_reg_9066_pp0_iter5_reg <= data_47_V_read_3_reg_9066_pp0_iter4_reg;
        data_47_V_read_3_reg_9066_pp0_iter6_reg <= data_47_V_read_3_reg_9066_pp0_iter5_reg;
        data_47_V_read_3_reg_9066_pp0_iter7_reg <= data_47_V_read_3_reg_9066_pp0_iter6_reg;
        data_47_V_read_3_reg_9066_pp0_iter8_reg <= data_47_V_read_3_reg_9066_pp0_iter7_reg;
        data_47_V_read_3_reg_9066_pp0_iter9_reg <= data_47_V_read_3_reg_9066_pp0_iter8_reg;
        data_48_V_read_3_reg_9040 <= data_48_V_read_int_reg;
        data_48_V_read_3_reg_9040_pp0_iter10_reg <= data_48_V_read_3_reg_9040_pp0_iter9_reg;
        data_48_V_read_3_reg_9040_pp0_iter11_reg <= data_48_V_read_3_reg_9040_pp0_iter10_reg;
        data_48_V_read_3_reg_9040_pp0_iter12_reg <= data_48_V_read_3_reg_9040_pp0_iter11_reg;
        data_48_V_read_3_reg_9040_pp0_iter13_reg <= data_48_V_read_3_reg_9040_pp0_iter12_reg;
        data_48_V_read_3_reg_9040_pp0_iter1_reg <= data_48_V_read_3_reg_9040;
        data_48_V_read_3_reg_9040_pp0_iter2_reg <= data_48_V_read_3_reg_9040_pp0_iter1_reg;
        data_48_V_read_3_reg_9040_pp0_iter3_reg <= data_48_V_read_3_reg_9040_pp0_iter2_reg;
        data_48_V_read_3_reg_9040_pp0_iter4_reg <= data_48_V_read_3_reg_9040_pp0_iter3_reg;
        data_48_V_read_3_reg_9040_pp0_iter5_reg <= data_48_V_read_3_reg_9040_pp0_iter4_reg;
        data_48_V_read_3_reg_9040_pp0_iter6_reg <= data_48_V_read_3_reg_9040_pp0_iter5_reg;
        data_48_V_read_3_reg_9040_pp0_iter7_reg <= data_48_V_read_3_reg_9040_pp0_iter6_reg;
        data_48_V_read_3_reg_9040_pp0_iter8_reg <= data_48_V_read_3_reg_9040_pp0_iter7_reg;
        data_48_V_read_3_reg_9040_pp0_iter9_reg <= data_48_V_read_3_reg_9040_pp0_iter8_reg;
        data_49_V_read_3_reg_9012 <= data_49_V_read_int_reg;
        data_49_V_read_3_reg_9012_pp0_iter10_reg <= data_49_V_read_3_reg_9012_pp0_iter9_reg;
        data_49_V_read_3_reg_9012_pp0_iter11_reg <= data_49_V_read_3_reg_9012_pp0_iter10_reg;
        data_49_V_read_3_reg_9012_pp0_iter12_reg <= data_49_V_read_3_reg_9012_pp0_iter11_reg;
        data_49_V_read_3_reg_9012_pp0_iter13_reg <= data_49_V_read_3_reg_9012_pp0_iter12_reg;
        data_49_V_read_3_reg_9012_pp0_iter1_reg <= data_49_V_read_3_reg_9012;
        data_49_V_read_3_reg_9012_pp0_iter2_reg <= data_49_V_read_3_reg_9012_pp0_iter1_reg;
        data_49_V_read_3_reg_9012_pp0_iter3_reg <= data_49_V_read_3_reg_9012_pp0_iter2_reg;
        data_49_V_read_3_reg_9012_pp0_iter4_reg <= data_49_V_read_3_reg_9012_pp0_iter3_reg;
        data_49_V_read_3_reg_9012_pp0_iter5_reg <= data_49_V_read_3_reg_9012_pp0_iter4_reg;
        data_49_V_read_3_reg_9012_pp0_iter6_reg <= data_49_V_read_3_reg_9012_pp0_iter5_reg;
        data_49_V_read_3_reg_9012_pp0_iter7_reg <= data_49_V_read_3_reg_9012_pp0_iter6_reg;
        data_49_V_read_3_reg_9012_pp0_iter8_reg <= data_49_V_read_3_reg_9012_pp0_iter7_reg;
        data_49_V_read_3_reg_9012_pp0_iter9_reg <= data_49_V_read_3_reg_9012_pp0_iter8_reg;
        data_4_V_read_10_reg_10273 <= data_4_V_read_int_reg;
        data_4_V_read_10_reg_10273_pp0_iter1_reg <= data_4_V_read_10_reg_10273;
        data_4_V_read_10_reg_10273_pp0_iter2_reg <= data_4_V_read_10_reg_10273_pp0_iter1_reg;
        data_4_V_read_10_reg_10273_pp0_iter3_reg <= data_4_V_read_10_reg_10273_pp0_iter2_reg;
        data_50_V_read51_reg_8984 <= data_50_V_read_int_reg;
        data_50_V_read51_reg_8984_pp0_iter10_reg <= data_50_V_read51_reg_8984_pp0_iter9_reg;
        data_50_V_read51_reg_8984_pp0_iter11_reg <= data_50_V_read51_reg_8984_pp0_iter10_reg;
        data_50_V_read51_reg_8984_pp0_iter12_reg <= data_50_V_read51_reg_8984_pp0_iter11_reg;
        data_50_V_read51_reg_8984_pp0_iter13_reg <= data_50_V_read51_reg_8984_pp0_iter12_reg;
        data_50_V_read51_reg_8984_pp0_iter14_reg <= data_50_V_read51_reg_8984_pp0_iter13_reg;
        data_50_V_read51_reg_8984_pp0_iter1_reg <= data_50_V_read51_reg_8984;
        data_50_V_read51_reg_8984_pp0_iter2_reg <= data_50_V_read51_reg_8984_pp0_iter1_reg;
        data_50_V_read51_reg_8984_pp0_iter3_reg <= data_50_V_read51_reg_8984_pp0_iter2_reg;
        data_50_V_read51_reg_8984_pp0_iter4_reg <= data_50_V_read51_reg_8984_pp0_iter3_reg;
        data_50_V_read51_reg_8984_pp0_iter5_reg <= data_50_V_read51_reg_8984_pp0_iter4_reg;
        data_50_V_read51_reg_8984_pp0_iter6_reg <= data_50_V_read51_reg_8984_pp0_iter5_reg;
        data_50_V_read51_reg_8984_pp0_iter7_reg <= data_50_V_read51_reg_8984_pp0_iter6_reg;
        data_50_V_read51_reg_8984_pp0_iter8_reg <= data_50_V_read51_reg_8984_pp0_iter7_reg;
        data_50_V_read51_reg_8984_pp0_iter9_reg <= data_50_V_read51_reg_8984_pp0_iter8_reg;
        data_51_V_read52_reg_8956 <= data_51_V_read_int_reg;
        data_51_V_read52_reg_8956_pp0_iter10_reg <= data_51_V_read52_reg_8956_pp0_iter9_reg;
        data_51_V_read52_reg_8956_pp0_iter11_reg <= data_51_V_read52_reg_8956_pp0_iter10_reg;
        data_51_V_read52_reg_8956_pp0_iter12_reg <= data_51_V_read52_reg_8956_pp0_iter11_reg;
        data_51_V_read52_reg_8956_pp0_iter13_reg <= data_51_V_read52_reg_8956_pp0_iter12_reg;
        data_51_V_read52_reg_8956_pp0_iter14_reg <= data_51_V_read52_reg_8956_pp0_iter13_reg;
        data_51_V_read52_reg_8956_pp0_iter1_reg <= data_51_V_read52_reg_8956;
        data_51_V_read52_reg_8956_pp0_iter2_reg <= data_51_V_read52_reg_8956_pp0_iter1_reg;
        data_51_V_read52_reg_8956_pp0_iter3_reg <= data_51_V_read52_reg_8956_pp0_iter2_reg;
        data_51_V_read52_reg_8956_pp0_iter4_reg <= data_51_V_read52_reg_8956_pp0_iter3_reg;
        data_51_V_read52_reg_8956_pp0_iter5_reg <= data_51_V_read52_reg_8956_pp0_iter4_reg;
        data_51_V_read52_reg_8956_pp0_iter6_reg <= data_51_V_read52_reg_8956_pp0_iter5_reg;
        data_51_V_read52_reg_8956_pp0_iter7_reg <= data_51_V_read52_reg_8956_pp0_iter6_reg;
        data_51_V_read52_reg_8956_pp0_iter8_reg <= data_51_V_read52_reg_8956_pp0_iter7_reg;
        data_51_V_read52_reg_8956_pp0_iter9_reg <= data_51_V_read52_reg_8956_pp0_iter8_reg;
        data_52_V_read_3_reg_8928 <= data_52_V_read_int_reg;
        data_52_V_read_3_reg_8928_pp0_iter10_reg <= data_52_V_read_3_reg_8928_pp0_iter9_reg;
        data_52_V_read_3_reg_8928_pp0_iter11_reg <= data_52_V_read_3_reg_8928_pp0_iter10_reg;
        data_52_V_read_3_reg_8928_pp0_iter12_reg <= data_52_V_read_3_reg_8928_pp0_iter11_reg;
        data_52_V_read_3_reg_8928_pp0_iter13_reg <= data_52_V_read_3_reg_8928_pp0_iter12_reg;
        data_52_V_read_3_reg_8928_pp0_iter14_reg <= data_52_V_read_3_reg_8928_pp0_iter13_reg;
        data_52_V_read_3_reg_8928_pp0_iter1_reg <= data_52_V_read_3_reg_8928;
        data_52_V_read_3_reg_8928_pp0_iter2_reg <= data_52_V_read_3_reg_8928_pp0_iter1_reg;
        data_52_V_read_3_reg_8928_pp0_iter3_reg <= data_52_V_read_3_reg_8928_pp0_iter2_reg;
        data_52_V_read_3_reg_8928_pp0_iter4_reg <= data_52_V_read_3_reg_8928_pp0_iter3_reg;
        data_52_V_read_3_reg_8928_pp0_iter5_reg <= data_52_V_read_3_reg_8928_pp0_iter4_reg;
        data_52_V_read_3_reg_8928_pp0_iter6_reg <= data_52_V_read_3_reg_8928_pp0_iter5_reg;
        data_52_V_read_3_reg_8928_pp0_iter7_reg <= data_52_V_read_3_reg_8928_pp0_iter6_reg;
        data_52_V_read_3_reg_8928_pp0_iter8_reg <= data_52_V_read_3_reg_8928_pp0_iter7_reg;
        data_52_V_read_3_reg_8928_pp0_iter9_reg <= data_52_V_read_3_reg_8928_pp0_iter8_reg;
        data_53_V_read_3_reg_8899 <= data_53_V_read_int_reg;
        data_53_V_read_3_reg_8899_pp0_iter10_reg <= data_53_V_read_3_reg_8899_pp0_iter9_reg;
        data_53_V_read_3_reg_8899_pp0_iter11_reg <= data_53_V_read_3_reg_8899_pp0_iter10_reg;
        data_53_V_read_3_reg_8899_pp0_iter12_reg <= data_53_V_read_3_reg_8899_pp0_iter11_reg;
        data_53_V_read_3_reg_8899_pp0_iter13_reg <= data_53_V_read_3_reg_8899_pp0_iter12_reg;
        data_53_V_read_3_reg_8899_pp0_iter14_reg <= data_53_V_read_3_reg_8899_pp0_iter13_reg;
        data_53_V_read_3_reg_8899_pp0_iter1_reg <= data_53_V_read_3_reg_8899;
        data_53_V_read_3_reg_8899_pp0_iter2_reg <= data_53_V_read_3_reg_8899_pp0_iter1_reg;
        data_53_V_read_3_reg_8899_pp0_iter3_reg <= data_53_V_read_3_reg_8899_pp0_iter2_reg;
        data_53_V_read_3_reg_8899_pp0_iter4_reg <= data_53_V_read_3_reg_8899_pp0_iter3_reg;
        data_53_V_read_3_reg_8899_pp0_iter5_reg <= data_53_V_read_3_reg_8899_pp0_iter4_reg;
        data_53_V_read_3_reg_8899_pp0_iter6_reg <= data_53_V_read_3_reg_8899_pp0_iter5_reg;
        data_53_V_read_3_reg_8899_pp0_iter7_reg <= data_53_V_read_3_reg_8899_pp0_iter6_reg;
        data_53_V_read_3_reg_8899_pp0_iter8_reg <= data_53_V_read_3_reg_8899_pp0_iter7_reg;
        data_53_V_read_3_reg_8899_pp0_iter9_reg <= data_53_V_read_3_reg_8899_pp0_iter8_reg;
        data_54_V_read_3_reg_8873 <= data_54_V_read_int_reg;
        data_54_V_read_3_reg_8873_pp0_iter10_reg <= data_54_V_read_3_reg_8873_pp0_iter9_reg;
        data_54_V_read_3_reg_8873_pp0_iter11_reg <= data_54_V_read_3_reg_8873_pp0_iter10_reg;
        data_54_V_read_3_reg_8873_pp0_iter12_reg <= data_54_V_read_3_reg_8873_pp0_iter11_reg;
        data_54_V_read_3_reg_8873_pp0_iter13_reg <= data_54_V_read_3_reg_8873_pp0_iter12_reg;
        data_54_V_read_3_reg_8873_pp0_iter14_reg <= data_54_V_read_3_reg_8873_pp0_iter13_reg;
        data_54_V_read_3_reg_8873_pp0_iter1_reg <= data_54_V_read_3_reg_8873;
        data_54_V_read_3_reg_8873_pp0_iter2_reg <= data_54_V_read_3_reg_8873_pp0_iter1_reg;
        data_54_V_read_3_reg_8873_pp0_iter3_reg <= data_54_V_read_3_reg_8873_pp0_iter2_reg;
        data_54_V_read_3_reg_8873_pp0_iter4_reg <= data_54_V_read_3_reg_8873_pp0_iter3_reg;
        data_54_V_read_3_reg_8873_pp0_iter5_reg <= data_54_V_read_3_reg_8873_pp0_iter4_reg;
        data_54_V_read_3_reg_8873_pp0_iter6_reg <= data_54_V_read_3_reg_8873_pp0_iter5_reg;
        data_54_V_read_3_reg_8873_pp0_iter7_reg <= data_54_V_read_3_reg_8873_pp0_iter6_reg;
        data_54_V_read_3_reg_8873_pp0_iter8_reg <= data_54_V_read_3_reg_8873_pp0_iter7_reg;
        data_54_V_read_3_reg_8873_pp0_iter9_reg <= data_54_V_read_3_reg_8873_pp0_iter8_reg;
        data_55_V_read_3_reg_8844 <= data_55_V_read_int_reg;
        data_55_V_read_3_reg_8844_pp0_iter10_reg <= data_55_V_read_3_reg_8844_pp0_iter9_reg;
        data_55_V_read_3_reg_8844_pp0_iter11_reg <= data_55_V_read_3_reg_8844_pp0_iter10_reg;
        data_55_V_read_3_reg_8844_pp0_iter12_reg <= data_55_V_read_3_reg_8844_pp0_iter11_reg;
        data_55_V_read_3_reg_8844_pp0_iter13_reg <= data_55_V_read_3_reg_8844_pp0_iter12_reg;
        data_55_V_read_3_reg_8844_pp0_iter14_reg <= data_55_V_read_3_reg_8844_pp0_iter13_reg;
        data_55_V_read_3_reg_8844_pp0_iter15_reg <= data_55_V_read_3_reg_8844_pp0_iter14_reg;
        data_55_V_read_3_reg_8844_pp0_iter1_reg <= data_55_V_read_3_reg_8844;
        data_55_V_read_3_reg_8844_pp0_iter2_reg <= data_55_V_read_3_reg_8844_pp0_iter1_reg;
        data_55_V_read_3_reg_8844_pp0_iter3_reg <= data_55_V_read_3_reg_8844_pp0_iter2_reg;
        data_55_V_read_3_reg_8844_pp0_iter4_reg <= data_55_V_read_3_reg_8844_pp0_iter3_reg;
        data_55_V_read_3_reg_8844_pp0_iter5_reg <= data_55_V_read_3_reg_8844_pp0_iter4_reg;
        data_55_V_read_3_reg_8844_pp0_iter6_reg <= data_55_V_read_3_reg_8844_pp0_iter5_reg;
        data_55_V_read_3_reg_8844_pp0_iter7_reg <= data_55_V_read_3_reg_8844_pp0_iter6_reg;
        data_55_V_read_3_reg_8844_pp0_iter8_reg <= data_55_V_read_3_reg_8844_pp0_iter7_reg;
        data_55_V_read_3_reg_8844_pp0_iter9_reg <= data_55_V_read_3_reg_8844_pp0_iter8_reg;
        data_56_V_read_3_reg_8814 <= data_56_V_read_int_reg;
        data_56_V_read_3_reg_8814_pp0_iter10_reg <= data_56_V_read_3_reg_8814_pp0_iter9_reg;
        data_56_V_read_3_reg_8814_pp0_iter11_reg <= data_56_V_read_3_reg_8814_pp0_iter10_reg;
        data_56_V_read_3_reg_8814_pp0_iter12_reg <= data_56_V_read_3_reg_8814_pp0_iter11_reg;
        data_56_V_read_3_reg_8814_pp0_iter13_reg <= data_56_V_read_3_reg_8814_pp0_iter12_reg;
        data_56_V_read_3_reg_8814_pp0_iter14_reg <= data_56_V_read_3_reg_8814_pp0_iter13_reg;
        data_56_V_read_3_reg_8814_pp0_iter15_reg <= data_56_V_read_3_reg_8814_pp0_iter14_reg;
        data_56_V_read_3_reg_8814_pp0_iter1_reg <= data_56_V_read_3_reg_8814;
        data_56_V_read_3_reg_8814_pp0_iter2_reg <= data_56_V_read_3_reg_8814_pp0_iter1_reg;
        data_56_V_read_3_reg_8814_pp0_iter3_reg <= data_56_V_read_3_reg_8814_pp0_iter2_reg;
        data_56_V_read_3_reg_8814_pp0_iter4_reg <= data_56_V_read_3_reg_8814_pp0_iter3_reg;
        data_56_V_read_3_reg_8814_pp0_iter5_reg <= data_56_V_read_3_reg_8814_pp0_iter4_reg;
        data_56_V_read_3_reg_8814_pp0_iter6_reg <= data_56_V_read_3_reg_8814_pp0_iter5_reg;
        data_56_V_read_3_reg_8814_pp0_iter7_reg <= data_56_V_read_3_reg_8814_pp0_iter6_reg;
        data_56_V_read_3_reg_8814_pp0_iter8_reg <= data_56_V_read_3_reg_8814_pp0_iter7_reg;
        data_56_V_read_3_reg_8814_pp0_iter9_reg <= data_56_V_read_3_reg_8814_pp0_iter8_reg;
        data_57_V_read_3_reg_8786 <= data_57_V_read_int_reg;
        data_57_V_read_3_reg_8786_pp0_iter10_reg <= data_57_V_read_3_reg_8786_pp0_iter9_reg;
        data_57_V_read_3_reg_8786_pp0_iter11_reg <= data_57_V_read_3_reg_8786_pp0_iter10_reg;
        data_57_V_read_3_reg_8786_pp0_iter12_reg <= data_57_V_read_3_reg_8786_pp0_iter11_reg;
        data_57_V_read_3_reg_8786_pp0_iter13_reg <= data_57_V_read_3_reg_8786_pp0_iter12_reg;
        data_57_V_read_3_reg_8786_pp0_iter14_reg <= data_57_V_read_3_reg_8786_pp0_iter13_reg;
        data_57_V_read_3_reg_8786_pp0_iter15_reg <= data_57_V_read_3_reg_8786_pp0_iter14_reg;
        data_57_V_read_3_reg_8786_pp0_iter1_reg <= data_57_V_read_3_reg_8786;
        data_57_V_read_3_reg_8786_pp0_iter2_reg <= data_57_V_read_3_reg_8786_pp0_iter1_reg;
        data_57_V_read_3_reg_8786_pp0_iter3_reg <= data_57_V_read_3_reg_8786_pp0_iter2_reg;
        data_57_V_read_3_reg_8786_pp0_iter4_reg <= data_57_V_read_3_reg_8786_pp0_iter3_reg;
        data_57_V_read_3_reg_8786_pp0_iter5_reg <= data_57_V_read_3_reg_8786_pp0_iter4_reg;
        data_57_V_read_3_reg_8786_pp0_iter6_reg <= data_57_V_read_3_reg_8786_pp0_iter5_reg;
        data_57_V_read_3_reg_8786_pp0_iter7_reg <= data_57_V_read_3_reg_8786_pp0_iter6_reg;
        data_57_V_read_3_reg_8786_pp0_iter8_reg <= data_57_V_read_3_reg_8786_pp0_iter7_reg;
        data_57_V_read_3_reg_8786_pp0_iter9_reg <= data_57_V_read_3_reg_8786_pp0_iter8_reg;
        data_58_V_read_3_reg_8756 <= data_58_V_read_int_reg;
        data_58_V_read_3_reg_8756_pp0_iter10_reg <= data_58_V_read_3_reg_8756_pp0_iter9_reg;
        data_58_V_read_3_reg_8756_pp0_iter11_reg <= data_58_V_read_3_reg_8756_pp0_iter10_reg;
        data_58_V_read_3_reg_8756_pp0_iter12_reg <= data_58_V_read_3_reg_8756_pp0_iter11_reg;
        data_58_V_read_3_reg_8756_pp0_iter13_reg <= data_58_V_read_3_reg_8756_pp0_iter12_reg;
        data_58_V_read_3_reg_8756_pp0_iter14_reg <= data_58_V_read_3_reg_8756_pp0_iter13_reg;
        data_58_V_read_3_reg_8756_pp0_iter15_reg <= data_58_V_read_3_reg_8756_pp0_iter14_reg;
        data_58_V_read_3_reg_8756_pp0_iter1_reg <= data_58_V_read_3_reg_8756;
        data_58_V_read_3_reg_8756_pp0_iter2_reg <= data_58_V_read_3_reg_8756_pp0_iter1_reg;
        data_58_V_read_3_reg_8756_pp0_iter3_reg <= data_58_V_read_3_reg_8756_pp0_iter2_reg;
        data_58_V_read_3_reg_8756_pp0_iter4_reg <= data_58_V_read_3_reg_8756_pp0_iter3_reg;
        data_58_V_read_3_reg_8756_pp0_iter5_reg <= data_58_V_read_3_reg_8756_pp0_iter4_reg;
        data_58_V_read_3_reg_8756_pp0_iter6_reg <= data_58_V_read_3_reg_8756_pp0_iter5_reg;
        data_58_V_read_3_reg_8756_pp0_iter7_reg <= data_58_V_read_3_reg_8756_pp0_iter6_reg;
        data_58_V_read_3_reg_8756_pp0_iter8_reg <= data_58_V_read_3_reg_8756_pp0_iter7_reg;
        data_58_V_read_3_reg_8756_pp0_iter9_reg <= data_58_V_read_3_reg_8756_pp0_iter8_reg;
        data_59_V_read_3_reg_8724 <= data_59_V_read_int_reg;
        data_59_V_read_3_reg_8724_pp0_iter10_reg <= data_59_V_read_3_reg_8724_pp0_iter9_reg;
        data_59_V_read_3_reg_8724_pp0_iter11_reg <= data_59_V_read_3_reg_8724_pp0_iter10_reg;
        data_59_V_read_3_reg_8724_pp0_iter12_reg <= data_59_V_read_3_reg_8724_pp0_iter11_reg;
        data_59_V_read_3_reg_8724_pp0_iter13_reg <= data_59_V_read_3_reg_8724_pp0_iter12_reg;
        data_59_V_read_3_reg_8724_pp0_iter14_reg <= data_59_V_read_3_reg_8724_pp0_iter13_reg;
        data_59_V_read_3_reg_8724_pp0_iter15_reg <= data_59_V_read_3_reg_8724_pp0_iter14_reg;
        data_59_V_read_3_reg_8724_pp0_iter16_reg <= data_59_V_read_3_reg_8724_pp0_iter15_reg;
        data_59_V_read_3_reg_8724_pp0_iter1_reg <= data_59_V_read_3_reg_8724;
        data_59_V_read_3_reg_8724_pp0_iter2_reg <= data_59_V_read_3_reg_8724_pp0_iter1_reg;
        data_59_V_read_3_reg_8724_pp0_iter3_reg <= data_59_V_read_3_reg_8724_pp0_iter2_reg;
        data_59_V_read_3_reg_8724_pp0_iter4_reg <= data_59_V_read_3_reg_8724_pp0_iter3_reg;
        data_59_V_read_3_reg_8724_pp0_iter5_reg <= data_59_V_read_3_reg_8724_pp0_iter4_reg;
        data_59_V_read_3_reg_8724_pp0_iter6_reg <= data_59_V_read_3_reg_8724_pp0_iter5_reg;
        data_59_V_read_3_reg_8724_pp0_iter7_reg <= data_59_V_read_3_reg_8724_pp0_iter6_reg;
        data_59_V_read_3_reg_8724_pp0_iter8_reg <= data_59_V_read_3_reg_8724_pp0_iter7_reg;
        data_59_V_read_3_reg_8724_pp0_iter9_reg <= data_59_V_read_3_reg_8724_pp0_iter8_reg;
        data_5_V_read_9_reg_10245 <= data_5_V_read_int_reg;
        data_5_V_read_9_reg_10245_pp0_iter1_reg <= data_5_V_read_9_reg_10245;
        data_5_V_read_9_reg_10245_pp0_iter2_reg <= data_5_V_read_9_reg_10245_pp0_iter1_reg;
        data_5_V_read_9_reg_10245_pp0_iter3_reg <= data_5_V_read_9_reg_10245_pp0_iter2_reg;
        data_60_V_read61_reg_8691 <= data_60_V_read_int_reg;
        data_60_V_read61_reg_8691_pp0_iter10_reg <= data_60_V_read61_reg_8691_pp0_iter9_reg;
        data_60_V_read61_reg_8691_pp0_iter11_reg <= data_60_V_read61_reg_8691_pp0_iter10_reg;
        data_60_V_read61_reg_8691_pp0_iter12_reg <= data_60_V_read61_reg_8691_pp0_iter11_reg;
        data_60_V_read61_reg_8691_pp0_iter13_reg <= data_60_V_read61_reg_8691_pp0_iter12_reg;
        data_60_V_read61_reg_8691_pp0_iter14_reg <= data_60_V_read61_reg_8691_pp0_iter13_reg;
        data_60_V_read61_reg_8691_pp0_iter15_reg <= data_60_V_read61_reg_8691_pp0_iter14_reg;
        data_60_V_read61_reg_8691_pp0_iter16_reg <= data_60_V_read61_reg_8691_pp0_iter15_reg;
        data_60_V_read61_reg_8691_pp0_iter1_reg <= data_60_V_read61_reg_8691;
        data_60_V_read61_reg_8691_pp0_iter2_reg <= data_60_V_read61_reg_8691_pp0_iter1_reg;
        data_60_V_read61_reg_8691_pp0_iter3_reg <= data_60_V_read61_reg_8691_pp0_iter2_reg;
        data_60_V_read61_reg_8691_pp0_iter4_reg <= data_60_V_read61_reg_8691_pp0_iter3_reg;
        data_60_V_read61_reg_8691_pp0_iter5_reg <= data_60_V_read61_reg_8691_pp0_iter4_reg;
        data_60_V_read61_reg_8691_pp0_iter6_reg <= data_60_V_read61_reg_8691_pp0_iter5_reg;
        data_60_V_read61_reg_8691_pp0_iter7_reg <= data_60_V_read61_reg_8691_pp0_iter6_reg;
        data_60_V_read61_reg_8691_pp0_iter8_reg <= data_60_V_read61_reg_8691_pp0_iter7_reg;
        data_60_V_read61_reg_8691_pp0_iter9_reg <= data_60_V_read61_reg_8691_pp0_iter8_reg;
        data_61_V_read62_reg_8663 <= data_61_V_read_int_reg;
        data_61_V_read62_reg_8663_pp0_iter10_reg <= data_61_V_read62_reg_8663_pp0_iter9_reg;
        data_61_V_read62_reg_8663_pp0_iter11_reg <= data_61_V_read62_reg_8663_pp0_iter10_reg;
        data_61_V_read62_reg_8663_pp0_iter12_reg <= data_61_V_read62_reg_8663_pp0_iter11_reg;
        data_61_V_read62_reg_8663_pp0_iter13_reg <= data_61_V_read62_reg_8663_pp0_iter12_reg;
        data_61_V_read62_reg_8663_pp0_iter14_reg <= data_61_V_read62_reg_8663_pp0_iter13_reg;
        data_61_V_read62_reg_8663_pp0_iter15_reg <= data_61_V_read62_reg_8663_pp0_iter14_reg;
        data_61_V_read62_reg_8663_pp0_iter16_reg <= data_61_V_read62_reg_8663_pp0_iter15_reg;
        data_61_V_read62_reg_8663_pp0_iter1_reg <= data_61_V_read62_reg_8663;
        data_61_V_read62_reg_8663_pp0_iter2_reg <= data_61_V_read62_reg_8663_pp0_iter1_reg;
        data_61_V_read62_reg_8663_pp0_iter3_reg <= data_61_V_read62_reg_8663_pp0_iter2_reg;
        data_61_V_read62_reg_8663_pp0_iter4_reg <= data_61_V_read62_reg_8663_pp0_iter3_reg;
        data_61_V_read62_reg_8663_pp0_iter5_reg <= data_61_V_read62_reg_8663_pp0_iter4_reg;
        data_61_V_read62_reg_8663_pp0_iter6_reg <= data_61_V_read62_reg_8663_pp0_iter5_reg;
        data_61_V_read62_reg_8663_pp0_iter7_reg <= data_61_V_read62_reg_8663_pp0_iter6_reg;
        data_61_V_read62_reg_8663_pp0_iter8_reg <= data_61_V_read62_reg_8663_pp0_iter7_reg;
        data_61_V_read62_reg_8663_pp0_iter9_reg <= data_61_V_read62_reg_8663_pp0_iter8_reg;
        data_62_V_read_3_reg_8645 <= data_62_V_read_int_reg;
        data_62_V_read_3_reg_8645_pp0_iter10_reg <= data_62_V_read_3_reg_8645_pp0_iter9_reg;
        data_62_V_read_3_reg_8645_pp0_iter11_reg <= data_62_V_read_3_reg_8645_pp0_iter10_reg;
        data_62_V_read_3_reg_8645_pp0_iter12_reg <= data_62_V_read_3_reg_8645_pp0_iter11_reg;
        data_62_V_read_3_reg_8645_pp0_iter13_reg <= data_62_V_read_3_reg_8645_pp0_iter12_reg;
        data_62_V_read_3_reg_8645_pp0_iter14_reg <= data_62_V_read_3_reg_8645_pp0_iter13_reg;
        data_62_V_read_3_reg_8645_pp0_iter15_reg <= data_62_V_read_3_reg_8645_pp0_iter14_reg;
        data_62_V_read_3_reg_8645_pp0_iter16_reg <= data_62_V_read_3_reg_8645_pp0_iter15_reg;
        data_62_V_read_3_reg_8645_pp0_iter1_reg <= data_62_V_read_3_reg_8645;
        data_62_V_read_3_reg_8645_pp0_iter2_reg <= data_62_V_read_3_reg_8645_pp0_iter1_reg;
        data_62_V_read_3_reg_8645_pp0_iter3_reg <= data_62_V_read_3_reg_8645_pp0_iter2_reg;
        data_62_V_read_3_reg_8645_pp0_iter4_reg <= data_62_V_read_3_reg_8645_pp0_iter3_reg;
        data_62_V_read_3_reg_8645_pp0_iter5_reg <= data_62_V_read_3_reg_8645_pp0_iter4_reg;
        data_62_V_read_3_reg_8645_pp0_iter6_reg <= data_62_V_read_3_reg_8645_pp0_iter5_reg;
        data_62_V_read_3_reg_8645_pp0_iter7_reg <= data_62_V_read_3_reg_8645_pp0_iter6_reg;
        data_62_V_read_3_reg_8645_pp0_iter8_reg <= data_62_V_read_3_reg_8645_pp0_iter7_reg;
        data_62_V_read_3_reg_8645_pp0_iter9_reg <= data_62_V_read_3_reg_8645_pp0_iter8_reg;
        data_63_V_read_3_reg_8620 <= data_63_V_read_int_reg;
        data_63_V_read_3_reg_8620_pp0_iter10_reg <= data_63_V_read_3_reg_8620_pp0_iter9_reg;
        data_63_V_read_3_reg_8620_pp0_iter11_reg <= data_63_V_read_3_reg_8620_pp0_iter10_reg;
        data_63_V_read_3_reg_8620_pp0_iter12_reg <= data_63_V_read_3_reg_8620_pp0_iter11_reg;
        data_63_V_read_3_reg_8620_pp0_iter13_reg <= data_63_V_read_3_reg_8620_pp0_iter12_reg;
        data_63_V_read_3_reg_8620_pp0_iter14_reg <= data_63_V_read_3_reg_8620_pp0_iter13_reg;
        data_63_V_read_3_reg_8620_pp0_iter15_reg <= data_63_V_read_3_reg_8620_pp0_iter14_reg;
        data_63_V_read_3_reg_8620_pp0_iter16_reg <= data_63_V_read_3_reg_8620_pp0_iter15_reg;
        data_63_V_read_3_reg_8620_pp0_iter1_reg <= data_63_V_read_3_reg_8620;
        data_63_V_read_3_reg_8620_pp0_iter2_reg <= data_63_V_read_3_reg_8620_pp0_iter1_reg;
        data_63_V_read_3_reg_8620_pp0_iter3_reg <= data_63_V_read_3_reg_8620_pp0_iter2_reg;
        data_63_V_read_3_reg_8620_pp0_iter4_reg <= data_63_V_read_3_reg_8620_pp0_iter3_reg;
        data_63_V_read_3_reg_8620_pp0_iter5_reg <= data_63_V_read_3_reg_8620_pp0_iter4_reg;
        data_63_V_read_3_reg_8620_pp0_iter6_reg <= data_63_V_read_3_reg_8620_pp0_iter5_reg;
        data_63_V_read_3_reg_8620_pp0_iter7_reg <= data_63_V_read_3_reg_8620_pp0_iter6_reg;
        data_63_V_read_3_reg_8620_pp0_iter8_reg <= data_63_V_read_3_reg_8620_pp0_iter7_reg;
        data_63_V_read_3_reg_8620_pp0_iter9_reg <= data_63_V_read_3_reg_8620_pp0_iter8_reg;
        data_6_V_read_9_reg_10218 <= data_6_V_read_int_reg;
        data_6_V_read_9_reg_10218_pp0_iter1_reg <= data_6_V_read_9_reg_10218;
        data_6_V_read_9_reg_10218_pp0_iter2_reg <= data_6_V_read_9_reg_10218_pp0_iter1_reg;
        data_6_V_read_9_reg_10218_pp0_iter3_reg <= data_6_V_read_9_reg_10218_pp0_iter2_reg;
        data_7_V_read_9_reg_10191 <= data_7_V_read_int_reg;
        data_7_V_read_9_reg_10191_pp0_iter1_reg <= data_7_V_read_9_reg_10191;
        data_7_V_read_9_reg_10191_pp0_iter2_reg <= data_7_V_read_9_reg_10191_pp0_iter1_reg;
        data_7_V_read_9_reg_10191_pp0_iter3_reg <= data_7_V_read_9_reg_10191_pp0_iter2_reg;
        data_7_V_read_9_reg_10191_pp0_iter4_reg <= data_7_V_read_9_reg_10191_pp0_iter3_reg;
        data_8_V_read_8_reg_10164 <= data_8_V_read_int_reg;
        data_8_V_read_8_reg_10164_pp0_iter1_reg <= data_8_V_read_8_reg_10164;
        data_8_V_read_8_reg_10164_pp0_iter2_reg <= data_8_V_read_8_reg_10164_pp0_iter1_reg;
        data_8_V_read_8_reg_10164_pp0_iter3_reg <= data_8_V_read_8_reg_10164_pp0_iter2_reg;
        data_8_V_read_8_reg_10164_pp0_iter4_reg <= data_8_V_read_8_reg_10164_pp0_iter3_reg;
        data_9_V_read_8_reg_10136 <= data_9_V_read_int_reg;
        data_9_V_read_8_reg_10136_pp0_iter1_reg <= data_9_V_read_8_reg_10136;
        data_9_V_read_8_reg_10136_pp0_iter2_reg <= data_9_V_read_8_reg_10136_pp0_iter1_reg;
        data_9_V_read_8_reg_10136_pp0_iter3_reg <= data_9_V_read_8_reg_10136_pp0_iter2_reg;
        data_9_V_read_8_reg_10136_pp0_iter4_reg <= data_9_V_read_8_reg_10136_pp0_iter3_reg;
        sub_ln703_106_reg_10707 <= sub_ln703_106_fu_1378_p2;
        sub_ln703_107_reg_10712 <= sub_ln703_107_fu_1383_p2;
        sub_ln703_108_reg_10717 <= sub_ln703_108_fu_1388_p2;
        sub_ln703_109_reg_10722 <= sub_ln703_109_fu_1407_p2;
        sub_ln703_10_reg_10420 <= sub_ln703_10_fu_615_p2;
        sub_ln703_115_reg_10727 <= sub_ln703_115_fu_1432_p2;
        sub_ln703_11_reg_10398 <= sub_ln703_11_fu_576_p2;
        sub_ln703_11_reg_10398_pp0_iter3_reg <= sub_ln703_11_reg_10398;
        sub_ln703_122_reg_10742 <= sub_ln703_122_fu_1462_p2;
        sub_ln703_123_reg_10747 <= sub_ln703_123_fu_1467_p2;
        sub_ln703_125_reg_10757 <= sub_ln703_125_fu_1482_p2;
        sub_ln703_128_reg_10762 <= sub_ln703_128_fu_1496_p2;
        sub_ln703_133_reg_10782 <= sub_ln703_133_fu_1532_p2;
        sub_ln703_137_reg_10787 <= sub_ln703_137_fu_1548_p2;
        sub_ln703_141_reg_10792 <= sub_ln703_141_fu_1553_p2;
        sub_ln703_142_reg_10797 <= sub_ln703_142_fu_1558_p2;
        sub_ln703_146_reg_10812 <= sub_ln703_146_fu_1580_p2;
        sub_ln703_152_reg_10822 <= sub_ln703_152_fu_1599_p2;
        sub_ln703_154_reg_10832 <= sub_ln703_154_fu_1609_p2;
        sub_ln703_15_reg_10430 <= sub_ln703_15_fu_631_p2;
        sub_ln703_166_reg_10863 <= sub_ln703_166_fu_1834_p2;
        sub_ln703_16_reg_10436 <= sub_ln703_16_fu_640_p2;
        sub_ln703_17_reg_10453 <= sub_ln703_17_fu_653_p2;
        sub_ln703_183_reg_10868 <= sub_ln703_183_fu_1959_p2;
        sub_ln703_184_reg_10878 <= sub_ln703_184_fu_1984_p2;
        sub_ln703_186_reg_10883 <= sub_ln703_186_fu_1994_p2;
        sub_ln703_18_reg_10459 <= sub_ln703_18_fu_658_p2;
        sub_ln703_191_reg_10893 <= sub_ln703_191_fu_2029_p2;
        sub_ln703_194_reg_10908 <= sub_ln703_194_fu_2054_p2;
        sub_ln703_196_reg_10913 <= sub_ln703_196_fu_2074_p2;
        sub_ln703_198_reg_10935 <= sub_ln703_198_fu_2099_p2;
        sub_ln703_1_reg_10348 <= sub_ln703_1_fu_540_p2;
        sub_ln703_200_reg_10950 <= sub_ln703_200_fu_2115_p2;
        sub_ln703_202_reg_10955 <= sub_ln703_202_fu_2120_p2;
        sub_ln703_203_reg_10965 <= sub_ln703_203_fu_2131_p2;
        sub_ln703_204_reg_10975 <= sub_ln703_204_fu_2142_p2;
        sub_ln703_208_reg_10985 <= sub_ln703_208_fu_2152_p2;
        sub_ln703_209_reg_10990 <= sub_ln703_209_fu_2157_p2;
        sub_ln703_20_reg_10465 <= sub_ln703_20_fu_662_p2;
        sub_ln703_210_reg_10995 <= sub_ln703_210_fu_2162_p2;
        sub_ln703_212_reg_11000 <= sub_ln703_212_fu_2173_p2;
        sub_ln703_230_reg_11010 <= sub_ln703_230_fu_2194_p2;
        sub_ln703_234_reg_11046 <= sub_ln703_234_fu_2395_p2;
        sub_ln703_237_reg_11020 <= sub_ln703_237_fu_2214_p2;
        sub_ln703_23_reg_10471 <= sub_ln703_23_fu_666_p2;
        sub_ln703_246_reg_11051 <= sub_ln703_246_fu_2477_p2;
        sub_ln703_249_reg_11056 <= sub_ln703_249_fu_2496_p2;
        sub_ln703_250_reg_11061 <= sub_ln703_250_fu_2501_p2;
        sub_ln703_251_reg_11066 <= sub_ln703_251_fu_2506_p2;
        sub_ln703_254_reg_11076 <= sub_ln703_254_fu_2525_p2;
        sub_ln703_256_reg_11081 <= sub_ln703_256_fu_2534_p2;
        sub_ln703_257_reg_11086 <= sub_ln703_257_fu_2539_p2;
        sub_ln703_261_reg_11091 <= sub_ln703_261_fu_2569_p2;
        sub_ln703_262_reg_11096 <= sub_ln703_262_fu_2574_p2;
        sub_ln703_263_reg_11101 <= sub_ln703_263_fu_2579_p2;
        sub_ln703_265_reg_11116 <= sub_ln703_265_fu_2613_p2;
        sub_ln703_270_reg_11121 <= sub_ln703_270_fu_2628_p2;
        sub_ln703_272_reg_11138 <= sub_ln703_272_fu_2647_p2;
        sub_ln703_274_reg_11143 <= sub_ln703_274_fu_2652_p2;
        sub_ln703_275_reg_11153 <= sub_ln703_275_fu_2662_p2;
        sub_ln703_281_reg_11163 <= sub_ln703_281_fu_2688_p2;
        sub_ln703_284_reg_11168 <= sub_ln703_284_fu_2698_p2;
        sub_ln703_289_reg_11173 <= sub_ln703_289_fu_2703_p2;
        sub_ln703_28_reg_10476 <= sub_ln703_28_fu_671_p2;
        sub_ln703_293_reg_11178 <= sub_ln703_293_fu_2708_p2;
        sub_ln703_296_reg_11183 <= sub_ln703_296_fu_2713_p2;
        sub_ln703_2_reg_10367 <= sub_ln703_2_fu_552_p2;
        sub_ln703_301_reg_11188 <= sub_ln703_301_fu_2718_p2;
        sub_ln703_313_reg_11257 <= sub_ln703_313_fu_2998_p2;
        sub_ln703_315_reg_11267 <= sub_ln703_315_fu_3021_p2;
        sub_ln703_326_reg_11277 <= sub_ln703_326_fu_3101_p2;
        sub_ln703_328_reg_11282 <= sub_ln703_328_fu_3111_p2;
        sub_ln703_333_reg_11292 <= sub_ln703_333_fu_3155_p2;
        sub_ln703_334_reg_11302 <= sub_ln703_334_fu_3175_p2;
        sub_ln703_336_reg_11307 <= sub_ln703_336_fu_3180_p2;
        sub_ln703_339_reg_11317 <= sub_ln703_339_fu_3200_p2;
        sub_ln703_340_reg_11322 <= sub_ln703_340_fu_3205_p2;
        sub_ln703_342_reg_11327 <= sub_ln703_342_fu_3215_p2;
        sub_ln703_344_reg_11332 <= sub_ln703_344_fu_3220_p2;
        sub_ln703_345_reg_11337 <= sub_ln703_345_fu_3234_p2;
        sub_ln703_350_reg_11342 <= sub_ln703_350_fu_3244_p2;
        sub_ln703_353_reg_11352 <= sub_ln703_353_fu_3269_p2;
        sub_ln703_356_reg_11367 <= sub_ln703_356_fu_3290_p2;
        sub_ln703_358_reg_11372 <= sub_ln703_358_fu_3300_p2;
        sub_ln703_362_reg_11377 <= sub_ln703_362_fu_3305_p2;
        sub_ln703_371_reg_11397 <= sub_ln703_371_fu_3324_p2;
        sub_ln703_384_reg_11474 <= sub_ln703_384_fu_3645_p2;
        sub_ln703_386_reg_11484 <= sub_ln703_386_fu_3660_p2;
        sub_ln703_387_reg_11489 <= sub_ln703_387_fu_3665_p2;
        sub_ln703_38_reg_10508 <= sub_ln703_38_fu_814_p2;
        sub_ln703_390_reg_11499 <= sub_ln703_390_fu_3690_p2;
        sub_ln703_393_reg_11504 <= sub_ln703_393_fu_3705_p2;
        sub_ln703_394_reg_11509 <= sub_ln703_394_fu_3710_p2;
        sub_ln703_395_reg_11514 <= sub_ln703_395_fu_3720_p2;
        sub_ln703_399_reg_11524 <= sub_ln703_399_fu_3761_p2;
        sub_ln703_39_reg_10513 <= sub_ln703_39_fu_819_p2;
        sub_ln703_3_reg_10379 <= sub_ln703_3_fu_560_p2;
        sub_ln703_401_reg_11529 <= sub_ln703_401_fu_3781_p2;
        sub_ln703_402_reg_11534 <= sub_ln703_402_fu_3786_p2;
        sub_ln703_403_reg_11539 <= sub_ln703_403_fu_3791_p2;
        sub_ln703_405_reg_11554 <= sub_ln703_405_fu_3816_p2;
        sub_ln703_408_reg_11564 <= sub_ln703_408_fu_3845_p2;
        sub_ln703_40_reg_10519 <= sub_ln703_40_fu_824_p2;
        sub_ln703_411_reg_11569 <= sub_ln703_411_fu_3850_p2;
        sub_ln703_412_reg_11574 <= sub_ln703_412_fu_3855_p2;
        sub_ln703_414_reg_11579 <= sub_ln703_414_fu_3860_p2;
        sub_ln703_416_reg_11584 <= sub_ln703_416_fu_3865_p2;
        sub_ln703_419_reg_11594 <= sub_ln703_419_fu_3884_p2;
        sub_ln703_43_reg_10524 <= sub_ln703_43_fu_838_p2;
        sub_ln703_440_reg_11624 <= sub_ln703_440_fu_3938_p2;
        sub_ln703_448_reg_11673 <= sub_ln703_448_fu_4206_p2;
        sub_ln703_452_reg_11678 <= sub_ln703_452_fu_4231_p2;
        sub_ln703_453_reg_11683 <= sub_ln703_453_fu_4236_p2;
        sub_ln703_458_reg_11688 <= sub_ln703_458_fu_4270_p2;
        sub_ln703_461_reg_11693 <= sub_ln703_461_fu_4303_p2;
        sub_ln703_462_reg_11703 <= sub_ln703_462_fu_4313_p2;
        sub_ln703_467_reg_11713 <= sub_ln703_467_fu_4333_p2;
        sub_ln703_468_reg_11718 <= sub_ln703_468_fu_4353_p2;
        sub_ln703_469_reg_11733 <= sub_ln703_469_fu_4368_p2;
        sub_ln703_470_reg_11738 <= sub_ln703_470_fu_4373_p2;
        sub_ln703_475_reg_11753 <= sub_ln703_475_fu_4418_p2;
        sub_ln703_482_reg_11773 <= sub_ln703_482_fu_4447_p2;
        sub_ln703_483_reg_11778 <= sub_ln703_483_fu_4452_p2;
        sub_ln703_488_reg_11783 <= sub_ln703_488_fu_4457_p2;
        sub_ln703_490_reg_11788 <= sub_ln703_490_fu_4462_p2;
        sub_ln703_491_reg_11793 <= sub_ln703_491_fu_4467_p2;
        sub_ln703_4_reg_10361 <= sub_ln703_4_fu_548_p2;
        sub_ln703_4_reg_10361_pp0_iter2_reg <= sub_ln703_4_reg_10361;
        sub_ln703_503_reg_11813 <= sub_ln703_503_fu_4516_p2;
        sub_ln703_505_reg_11818 <= sub_ln703_505_fu_4521_p2;
        sub_ln703_526_reg_11864 <= sub_ln703_526_fu_4860_p2;
        sub_ln703_527_reg_11869 <= sub_ln703_527_fu_4865_p2;
        sub_ln703_529_reg_11879 <= sub_ln703_529_fu_4880_p2;
        sub_ln703_532_reg_11884 <= sub_ln703_532_fu_4894_p2;
        sub_ln703_533_reg_11894 <= sub_ln703_533_fu_4904_p2;
        sub_ln703_535_reg_11899 <= sub_ln703_535_fu_4919_p2;
        sub_ln703_538_reg_11904 <= sub_ln703_538_fu_4934_p2;
        sub_ln703_539_reg_11909 <= sub_ln703_539_fu_4939_p2;
        sub_ln703_53_reg_10534 <= sub_ln703_53_fu_912_p2;
        sub_ln703_540_reg_11914 <= sub_ln703_540_fu_4944_p2;
        sub_ln703_541_reg_11919 <= sub_ln703_541_fu_4949_p2;
        sub_ln703_542_reg_11924 <= sub_ln703_542_fu_4954_p2;
        sub_ln703_544_reg_11934 <= sub_ln703_544_fu_4984_p2;
        sub_ln703_551_reg_11949 <= sub_ln703_551_fu_5004_p2;
        sub_ln703_556_reg_11964 <= sub_ln703_556_fu_5024_p2;
        sub_ln703_557_reg_11969 <= sub_ln703_557_fu_5029_p2;
        sub_ln703_558_reg_11974 <= sub_ln703_558_fu_5034_p2;
        sub_ln703_573_reg_12007 <= sub_ln703_573_fu_5101_p2;
        sub_ln703_582_reg_12012 <= sub_ln703_582_fu_5106_p2;
        sub_ln703_583_reg_12017 <= sub_ln703_583_fu_5111_p2;
        sub_ln703_586_reg_12061 <= sub_ln703_586_fu_5351_p2;
        sub_ln703_589_reg_12066 <= sub_ln703_589_fu_5375_p2;
        sub_ln703_58_reg_10545 <= sub_ln703_58_fu_922_p2;
        sub_ln703_593_reg_12071 <= sub_ln703_593_fu_5410_p2;
        sub_ln703_594_reg_12076 <= sub_ln703_594_fu_5415_p2;
        sub_ln703_595_reg_12081 <= sub_ln703_595_fu_5420_p2;
        sub_ln703_598_reg_12091 <= sub_ln703_598_fu_5454_p2;
        sub_ln703_603_reg_12101 <= sub_ln703_603_fu_5491_p2;
        sub_ln703_604_reg_12106 <= sub_ln703_604_fu_5496_p2;
        sub_ln703_605_reg_12111 <= sub_ln703_605_fu_5501_p2;
        sub_ln703_608_reg_12116 <= sub_ln703_608_fu_5511_p2;
        sub_ln703_609_reg_12121 <= sub_ln703_609_fu_5516_p2;
        sub_ln703_610_reg_12126 <= sub_ln703_610_fu_5521_p2;
        sub_ln703_612_reg_12131 <= sub_ln703_612_fu_5526_p2;
        sub_ln703_613_reg_12136 <= sub_ln703_613_fu_5531_p2;
        sub_ln703_614_reg_12141 <= sub_ln703_614_fu_5536_p2;
        sub_ln703_618_reg_12156 <= sub_ln703_618_fu_5566_p2;
        sub_ln703_624_reg_12166 <= sub_ln703_624_fu_5596_p2;
        sub_ln703_62_reg_10550 <= sub_ln703_62_fu_942_p2;
        sub_ln703_630_reg_12171 <= sub_ln703_630_fu_5627_p2;
        sub_ln703_631_reg_12176 <= sub_ln703_631_fu_5632_p2;
        sub_ln703_634_reg_12181 <= sub_ln703_634_fu_5637_p2;
        sub_ln703_637_reg_12186 <= sub_ln703_637_fu_5642_p2;
        sub_ln703_638_reg_12191 <= sub_ln703_638_fu_5647_p2;
        sub_ln703_63_reg_10555 <= sub_ln703_63_fu_947_p2;
        sub_ln703_644_reg_12204 <= sub_ln703_644_fu_5656_p2;
        sub_ln703_648_reg_12209 <= sub_ln703_648_fu_5661_p2;
        sub_ln703_64_reg_10560 <= sub_ln703_64_fu_957_p2;
        sub_ln703_650_reg_12214 <= sub_ln703_650_fu_5666_p2;
        sub_ln703_662_reg_12248 <= sub_ln703_662_fu_5918_p2;
        sub_ln703_665_reg_12253 <= sub_ln703_665_fu_5932_p2;
        sub_ln703_667_reg_12263 <= sub_ln703_667_fu_5956_p2;
        sub_ln703_669_reg_12268 <= sub_ln703_669_fu_5975_p2;
        sub_ln703_66_reg_10581 <= sub_ln703_66_fu_987_p2;
        sub_ln703_676_reg_12278 <= sub_ln703_676_fu_6033_p2;
        sub_ln703_678_reg_12283 <= sub_ln703_678_fu_6052_p2;
        sub_ln703_679_reg_12288 <= sub_ln703_679_fu_6057_p2;
        sub_ln703_680_reg_12293 <= sub_ln703_680_fu_6062_p2;
        sub_ln703_682_reg_12298 <= sub_ln703_682_fu_6067_p2;
        sub_ln703_684_reg_12303 <= sub_ln703_684_fu_6072_p2;
        sub_ln703_686_reg_12308 <= sub_ln703_686_fu_6077_p2;
        sub_ln703_687_reg_12313 <= sub_ln703_687_fu_6086_p2;
        sub_ln703_688_reg_12318 <= sub_ln703_688_fu_6091_p2;
        sub_ln703_690_reg_12323 <= sub_ln703_690_fu_6101_p2;
        sub_ln703_691_reg_12328 <= sub_ln703_691_fu_6106_p2;
        sub_ln703_692_reg_12333 <= sub_ln703_692_fu_6111_p2;
        sub_ln703_693_reg_12338 <= sub_ln703_693_fu_6116_p2;
        sub_ln703_694_reg_12343 <= sub_ln703_694_fu_6126_p2;
        sub_ln703_696_reg_12353 <= sub_ln703_696_fu_6136_p2;
        sub_ln703_697_reg_12358 <= sub_ln703_697_fu_6141_p2;
        sub_ln703_6_reg_10408 <= sub_ln703_6_fu_595_p2;
        sub_ln703_700_reg_12378 <= sub_ln703_700_fu_6172_p2;
        sub_ln703_704_reg_12383 <= sub_ln703_704_fu_6177_p2;
        sub_ln703_707_reg_12388 <= sub_ln703_707_fu_6182_p2;
        sub_ln703_70_reg_10586 <= sub_ln703_70_fu_992_p2;
        sub_ln703_71_reg_10596 <= sub_ln703_71_fu_1002_p2;
        sub_ln703_724_reg_12450 <= sub_ln703_724_fu_6432_p2;
        sub_ln703_727_reg_12460 <= sub_ln703_727_fu_6452_p2;
        sub_ln703_728_reg_12465 <= sub_ln703_728_fu_6457_p2;
        sub_ln703_733_reg_12470 <= sub_ln703_733_fu_6487_p2;
        sub_ln703_736_reg_12475 <= sub_ln703_736_fu_6502_p2;
        sub_ln703_73_reg_10611 <= sub_ln703_73_fu_1026_p2;
        sub_ln703_746_reg_12500 <= sub_ln703_746_fu_6579_p2;
        sub_ln703_749_reg_12510 <= sub_ln703_749_fu_6599_p2;
        sub_ln703_757_reg_12515 <= sub_ln703_757_fu_6629_p2;
        sub_ln703_759_reg_12525 <= sub_ln703_759_fu_6639_p2;
        sub_ln703_75_reg_10616 <= sub_ln703_75_fu_1031_p2;
        sub_ln703_761_reg_12530 <= sub_ln703_761_fu_6644_p2;
        sub_ln703_763_reg_12540 <= sub_ln703_763_fu_6654_p2;
        sub_ln703_767_reg_12545 <= sub_ln703_767_fu_6659_p2;
        sub_ln703_769_reg_12555 <= sub_ln703_769_fu_6684_p2;
        sub_ln703_770_reg_12570 <= sub_ln703_770_fu_6708_p2;
        sub_ln703_781_reg_12580 <= sub_ln703_781_fu_6739_p2;
        sub_ln703_787_reg_12590 <= sub_ln703_787_fu_6759_p2;
        sub_ln703_797_reg_12645 <= sub_ln703_797_fu_7030_p2;
        sub_ln703_799_reg_12595 <= sub_ln703_799_fu_6764_p2;
        sub_ln703_801_reg_12660 <= sub_ln703_801_fu_7060_p2;
        sub_ln703_802_reg_12665 <= sub_ln703_802_fu_7065_p2;
        sub_ln703_805_reg_12670 <= sub_ln703_805_fu_7079_p2;
        sub_ln703_807_reg_12685 <= sub_ln703_807_fu_7099_p2;
        sub_ln703_808_reg_12700 <= sub_ln703_808_fu_7137_p2;
        sub_ln703_814_reg_12735 <= sub_ln703_814_fu_7200_p2;
        sub_ln703_816_reg_12740 <= sub_ln703_816_fu_7205_p2;
        sub_ln703_818_reg_12745 <= sub_ln703_818_fu_7210_p2;
        sub_ln703_820_reg_12750 <= sub_ln703_820_fu_7215_p2;
        sub_ln703_821_reg_12755 <= sub_ln703_821_fu_7220_p2;
        sub_ln703_823_reg_12760 <= sub_ln703_823_fu_7225_p2;
        sub_ln703_824_reg_12765 <= sub_ln703_824_fu_7230_p2;
        sub_ln703_825_reg_12770 <= sub_ln703_825_fu_7235_p2;
        sub_ln703_852_reg_12790 <= sub_ln703_852_fu_7319_p2;
        sub_ln703_857_reg_12835 <= sub_ln703_857_fu_7600_p2;
        sub_ln703_858_reg_12840 <= sub_ln703_858_fu_7605_p2;
        sub_ln703_859_reg_12850 <= sub_ln703_859_fu_7615_p2;
        sub_ln703_862_reg_12795 <= sub_ln703_862_fu_7324_p2;
        sub_ln703_863_reg_12860 <= sub_ln703_863_fu_7639_p2;
        sub_ln703_865_reg_12865 <= sub_ln703_865_fu_7649_p2;
        sub_ln703_866_reg_12870 <= sub_ln703_866_fu_7654_p2;
        sub_ln703_867_reg_12880 <= sub_ln703_867_fu_7669_p2;
        sub_ln703_868_reg_12885 <= sub_ln703_868_fu_7674_p2;
        sub_ln703_869_reg_12800 <= sub_ln703_869_fu_7329_p2;
        sub_ln703_869_reg_12800_pp0_iter16_reg <= sub_ln703_869_reg_12800;
        sub_ln703_870_reg_12895 <= sub_ln703_870_fu_7685_p2;
        sub_ln703_873_reg_12900 <= sub_ln703_873_fu_7710_p2;
        sub_ln703_875_reg_12910 <= sub_ln703_875_fu_7730_p2;
        sub_ln703_879_reg_12915 <= sub_ln703_879_fu_7735_p2;
        sub_ln703_880_reg_12920 <= sub_ln703_880_fu_7750_p2;
        sub_ln703_881_reg_12925 <= sub_ln703_881_fu_7755_p2;
        sub_ln703_892_reg_12935 <= sub_ln703_892_fu_7780_p2;
        sub_ln703_893_reg_12940 <= sub_ln703_893_fu_7785_p2;
        sub_ln703_894_reg_12945 <= sub_ln703_894_fu_7790_p2;
        sub_ln703_895_reg_12950 <= sub_ln703_895_fu_7795_p2;
        sub_ln703_898_reg_12955 <= sub_ln703_898_fu_7805_p2;
        sub_ln703_8_reg_10392 <= sub_ln703_8_fu_572_p2;
        sub_ln703_904_reg_12960 <= sub_ln703_904_fu_7810_p2;
        sub_ln703_911_reg_12970 <= sub_ln703_911_fu_7833_p2;
        sub_ln703_917_reg_12975 <= sub_ln703_917_fu_7838_p2;
        sub_ln703_922_reg_12980 <= sub_ln703_922_fu_7843_p2;
        sub_ln703_92_reg_10636 <= sub_ln703_92_fu_1054_p2;
        sub_ln703_96_reg_10677 <= sub_ln703_96_fu_1294_p2;
        sub_ln703_98_reg_10697 <= sub_ln703_98_fu_1319_p2;
        sub_ln703_reg_10342 <= sub_ln703_fu_536_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_986_fu_8255_p2;
        ap_return_10_int_reg <= acc_10_V_fu_8310_p2;
        ap_return_11_int_reg <= acc_11_V_fu_8315_p2;
        ap_return_12_int_reg <= acc_12_V_fu_8320_p2;
        ap_return_13_int_reg <= acc_13_V_fu_8330_p2;
        ap_return_14_int_reg <= acc_14_V_fu_8335_p2;
        ap_return_15_int_reg <= acc_15_V_fu_8340_p2;
        ap_return_16_int_reg <= acc_16_V_fu_8345_p2;
        ap_return_17_int_reg <= acc_17_V_fu_8350_p2;
        ap_return_18_int_reg <= acc_18_V_fu_8355_p2;
        ap_return_19_int_reg <= acc_19_V_fu_8360_p2;
        ap_return_1_int_reg <= acc_1_V_fu_8265_p2;
        ap_return_20_int_reg <= acc_20_V_fu_8365_p2;
        ap_return_21_int_reg <= acc_21_V_reg_12991;
        ap_return_22_int_reg <= acc_22_V_fu_8370_p2;
        ap_return_23_int_reg <= acc_23_V_fu_8375_p2;
        ap_return_24_int_reg <= acc_24_V_fu_8380_p2;
        ap_return_25_int_reg <= acc_25_V_fu_8385_p2;
        ap_return_26_int_reg <= acc_26_V_fu_8390_p2;
        ap_return_27_int_reg <= acc_27_V_fu_8400_p2;
        ap_return_28_int_reg <= acc_28_V_fu_8405_p2;
        ap_return_29_int_reg <= acc_29_V_fu_8414_p2;
        ap_return_2_int_reg <= acc_2_V_fu_8270_p2;
        ap_return_30_int_reg <= acc_30_V_fu_8419_p2;
        ap_return_31_int_reg <= acc_31_V_fu_8424_p2;
        ap_return_3_int_reg <= acc_3_V_fu_8275_p2;
        ap_return_4_int_reg <= acc_4_V_fu_8280_p2;
        ap_return_5_int_reg <= acc_5_V_fu_8285_p2;
        ap_return_6_int_reg <= acc_6_V_fu_8290_p2;
        ap_return_7_int_reg <= acc_7_V_fu_8295_p2;
        ap_return_8_int_reg <= acc_8_V_fu_8300_p2;
        ap_return_9_int_reg <= acc_9_V_fu_8305_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_32_V_read_int_reg <= data_32_V_read;
        data_33_V_read_int_reg <= data_33_V_read;
        data_34_V_read_int_reg <= data_34_V_read;
        data_35_V_read_int_reg <= data_35_V_read;
        data_36_V_read_int_reg <= data_36_V_read;
        data_37_V_read_int_reg <= data_37_V_read;
        data_38_V_read_int_reg <= data_38_V_read;
        data_39_V_read_int_reg <= data_39_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_40_V_read_int_reg <= data_40_V_read;
        data_41_V_read_int_reg <= data_41_V_read;
        data_42_V_read_int_reg <= data_42_V_read;
        data_43_V_read_int_reg <= data_43_V_read;
        data_44_V_read_int_reg <= data_44_V_read;
        data_45_V_read_int_reg <= data_45_V_read;
        data_46_V_read_int_reg <= data_46_V_read;
        data_47_V_read_int_reg <= data_47_V_read;
        data_48_V_read_int_reg <= data_48_V_read;
        data_49_V_read_int_reg <= data_49_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_50_V_read_int_reg <= data_50_V_read;
        data_51_V_read_int_reg <= data_51_V_read;
        data_52_V_read_int_reg <= data_52_V_read;
        data_53_V_read_int_reg <= data_53_V_read;
        data_54_V_read_int_reg <= data_54_V_read;
        data_55_V_read_int_reg <= data_55_V_read;
        data_56_V_read_int_reg <= data_56_V_read;
        data_57_V_read_int_reg <= data_57_V_read;
        data_58_V_read_int_reg <= data_58_V_read;
        data_59_V_read_int_reg <= data_59_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_60_V_read_int_reg <= data_60_V_read;
        data_61_V_read_int_reg <= data_61_V_read;
        data_62_V_read_int_reg <= data_62_V_read;
        data_63_V_read_int_reg <= data_63_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_986_fu_8255_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_8265_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = acc_10_V_fu_8310_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = acc_11_V_fu_8315_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = acc_12_V_fu_8320_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = acc_13_V_fu_8330_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = acc_14_V_fu_8335_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = acc_15_V_fu_8340_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = acc_16_V_fu_8345_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = acc_17_V_fu_8350_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = acc_18_V_fu_8355_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = acc_19_V_fu_8360_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_8270_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = acc_20_V_fu_8365_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = acc_21_V_reg_12991;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = acc_22_V_fu_8370_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = acc_23_V_fu_8375_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = acc_24_V_fu_8380_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = acc_25_V_fu_8385_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = acc_26_V_fu_8390_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = acc_27_V_fu_8400_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = acc_28_V_fu_8405_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = acc_29_V_fu_8414_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_8275_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = acc_30_V_fu_8419_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = acc_31_V_fu_8424_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_8280_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = acc_5_V_fu_8285_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = acc_6_V_fu_8290_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = acc_7_V_fu_8295_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = acc_8_V_fu_8300_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = acc_9_V_fu_8305_p2;
    end
end

assign acc_10_V_fu_8310_p2 = (add_ln703_974_fu_8159_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_11_V_fu_8315_p2 = (sub_ln703_934_fu_8165_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_12_V_fu_8320_p2 = (add_ln703_976_fu_8175_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_13_V_fu_8330_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_994_fu_8325_p2);

assign acc_14_V_fu_8335_p2 = (sub_ln703_935_fu_8181_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_15_V_fu_8340_p2 = (add_ln703_978_fu_8191_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_16_V_fu_8345_p2 = (add_ln703_979_fu_8197_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_17_V_fu_8350_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_924_fu_8072_p2);

assign acc_18_V_fu_8355_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_925_fu_8076_p2);

assign acc_19_V_fu_8360_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_926_fu_8080_p2);

assign acc_1_V_fu_8265_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_987_fu_8260_p2);

assign acc_20_V_fu_8365_p2 = (add_ln703_980_fu_8203_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_21_V_fu_7872_p2 = (add_ln703_1003_fu_7867_p2 + add_ln703_1001_fu_7857_p2);

assign acc_22_V_fu_8370_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_927_fu_8085_p2);

assign acc_23_V_fu_8375_p2 = (sub_ln703_936_fu_8209_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_24_V_fu_8380_p2 = (add_ln703_981_fu_8214_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_25_V_fu_8385_p2 = (sub_ln703_937_fu_8219_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_26_V_fu_8390_p2 = (sub_ln703_938_fu_8224_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_27_V_fu_8400_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_1007_fu_8395_p2);

assign acc_28_V_fu_8405_p2 = (sub_ln703_939_fu_8229_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_29_V_fu_8414_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_1009_fu_8410_p2);

assign acc_2_V_fu_8270_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_919_fu_8037_p2);

assign acc_30_V_fu_8419_p2 = (sub_ln703_940_fu_8234_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_31_V_fu_8424_p2 = (add_ln703_983_fu_8244_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_3_V_fu_8275_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_920_fu_8042_p2);

assign acc_4_V_fu_8280_p2 = (sub_ln703_930_fu_8120_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_5_V_fu_8285_p2 = (add_ln703_971_fu_8129_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_6_V_fu_8290_p2 = (sub_ln703_931_fu_8134_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_7_V_fu_8295_p2 = (sub_ln703_932_fu_8139_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_8_V_fu_8300_p2 = (sub_ln703_933_fu_8143_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_9_V_fu_8305_p2 = (add_ln703_973_fu_8153_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign add_ln703_1000_fu_7852_p2 = (sub_ln703_819_fu_7386_p2 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_1001_fu_7857_p2 = (add_ln703_937_fu_7659_p2 + add_ln703_1000_fu_7852_p2);

assign add_ln703_1002_fu_7863_p2 = (add_ln703_985_reg_12819 + data_61_V_read62_reg_8663_pp0_iter15_reg);

assign add_ln703_1003_fu_7867_p2 = (add_ln703_1002_fu_7863_p2 + add_ln703_954_reg_12812);

assign add_ln703_1007_fu_8395_p2 = (sub_ln703_916_fu_8028_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_1009_fu_8410_p2 = (sub_ln703_917_reg_12975 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_130_fu_556_p2 = (sub_ln703_1_reg_10348 + data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign add_ln703_131_fu_544_p2 = (add_ln703_reg_10335 + data_2_V_read_10_reg_10312);

assign add_ln703_132_fu_599_p2 = (add_ln703_130_reg_10373 + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_133_fu_603_p2 = (sub_ln703_3_reg_10379 + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_134_fu_568_p2 = (add_ln703_131_reg_10354 + data_3_V_read_10_reg_10295_pp0_iter1_reg);

assign add_ln703_135_fu_619_p2 = (sub_ln703_2_reg_10367 + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_136_fu_623_p2 = (sub_ln703_4_reg_10361_pp0_iter2_reg + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_137_fu_697_p2 = (sub_ln703_6_reg_10408 + data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign add_ln703_138_fu_701_p2 = (add_ln703_132_reg_10414 + data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign add_ln703_139_fu_636_p2 = (add_ln703_134_reg_10385 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_140_fu_644_p2 = (sub_ln703_7_fu_607_p2 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_141_fu_649_p2 = (sub_ln703_8_reg_10392 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_142_fu_581_p2 = (sub_ln703_reg_10342 + data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign add_ln703_143_fu_585_p2 = (data_3_V_read_10_reg_10295_pp0_iter1_reg + data_4_V_read_10_reg_10273_pp0_iter1_reg);

assign add_ln703_144_fu_589_p2 = (add_ln703_143_fu_585_p2 + add_ln703_142_fu_581_p2);

assign add_ln703_145_fu_736_p2 = (add_ln703_138_fu_701_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_146_fu_741_p2 = (sub_ln703_15_reg_10430 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_147_fu_745_p2 = (sub_ln703_16_reg_10436 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_148_fu_757_p2 = (add_ln703_141_reg_10447 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_149_fu_773_p2 = (sub_ln703_19_fu_705_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_150_fu_782_p2 = (sub_ln703_22_fu_713_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_151_fu_791_p2 = (sub_ln703_20_reg_10465 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_152_fu_804_p2 = (sub_ln703_24_fu_717_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_153_fu_809_p2 = (sub_ln703_25_fu_722_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_154_fu_843_p2 = (sub_ln703_30_fu_753_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_155_fu_868_p2 = (data_5_V_read_9_reg_10245_pp0_iter3_reg + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_156_fu_872_p2 = (add_ln703_155_fu_868_p2 + sub_ln703_18_reg_10459);

assign add_ln703_157_fu_892_p2 = (sub_ln703_35_fu_787_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_158_fu_676_p2 = (sub_ln703_12_fu_627_p2 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_160_fu_902_p2 = (add_ln703_155_fu_868_p2 + add_ln703_158_reg_10482);

assign add_ln703_161_fu_681_p2 = (data_6_V_read_9_reg_10218_pp0_iter2_reg + data_7_V_read_9_reg_10191_pp0_iter2_reg);

assign add_ln703_162_fu_917_p2 = (add_ln703_161_reg_10487 + sub_ln703_26_fu_727_p2);

assign add_ln703_163_fu_1098_p2 = (sub_ln703_39_reg_10513 + data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign add_ln703_164_fu_937_p2 = (sub_ln703_45_fu_853_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_165_fu_952_p2 = (sub_ln703_38_fu_814_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_166_fu_962_p2 = (sub_ln703_21_fu_709_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_168_fu_967_p2 = (add_ln703_161_reg_10487 + add_ln703_166_fu_962_p2);

assign add_ln703_170_fu_972_p2 = (add_ln703_161_reg_10487 + add_ln703_149_fu_773_p2);

assign add_ln703_171_fu_977_p2 = (sub_ln703_51_fu_897_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_173_fu_982_p2 = (add_ln703_161_reg_10487 + sub_ln703_36_fu_795_p2);

assign add_ln703_174_fu_1114_p2 = (sub_ln703_54_fu_1086_p2 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_175_fu_1123_p2 = (sub_ln703_55_fu_1090_p2 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_176_fu_1128_p2 = (sub_ln703_56_fu_1094_p2 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_177_fu_997_p2 = (sub_ln703_61_fu_932_p2 + data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign add_ln703_178_fu_1007_p2 = (sub_ln703_17_reg_10453 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_179_fu_685_p2 = (data_7_V_read_9_reg_10191_pp0_iter2_reg + data_8_V_read_8_reg_10164_pp0_iter2_reg);

assign add_ln703_180_fu_1011_p2 = (add_ln703_179_reg_10495 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_181_fu_1015_p2 = (add_ln703_180_fu_1011_p2 + add_ln703_178_fu_1007_p2);

assign add_ln703_183_fu_1021_p2 = (add_ln703_179_reg_10495 + sub_ln703_47_fu_863_p2);

assign add_ln703_184_fu_1143_p2 = (sub_ln703_62_reg_10550 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_186_fu_1036_p2 = (add_ln703_179_reg_10495 + sub_ln703_50_fu_887_p2);

assign add_ln703_187_fu_1041_p2 = (sub_ln703_28_reg_10476 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_189_fu_1045_p2 = (add_ln703_179_reg_10495 + add_ln703_187_fu_1041_p2);

assign add_ln703_190_fu_1172_p2 = (sub_ln703_64_reg_10560 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_191_fu_1176_p2 = (sub_ln703_66_reg_10581 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_192_fu_1050_p2 = (data_8_V_read_8_reg_10164_pp0_iter3_reg + data_9_V_read_8_reg_10136_pp0_iter3_reg);

assign add_ln703_193_fu_1180_p2 = (add_ln703_192_reg_10626 + sub_ln703_53_reg_10534);

assign add_ln703_194_fu_1189_p2 = (sub_ln703_67_fu_1119_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_195_fu_1204_p2 = (sub_ln703_69_fu_1138_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_197_fu_1209_p2 = (add_ln703_192_reg_10626 + sub_ln703_58_reg_10545);

assign add_ln703_199_fu_1213_p2 = (add_ln703_192_reg_10626 + sub_ln703_59_fu_1106_p2);

assign add_ln703_200_fu_1226_p2 = (sub_ln703_71_reg_10596 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_201_fu_1243_p2 = (sub_ln703_72_fu_1147_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_202_fu_1265_p2 = (sub_ln703_77_fu_1159_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_203_fu_1270_p2 = (sub_ln703_78_fu_1164_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_204_fu_1059_p2 = (sub_ln703_52_fu_907_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_206_fu_1290_p2 = (add_ln703_192_reg_10626 + add_ln703_204_reg_10641);

assign add_ln703_207_fu_1299_p2 = (sub_ln703_80_fu_1184_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_208_fu_1309_p2 = (sub_ln703_82_fu_1199_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_209_fu_1064_p2 = (data_9_V_read_8_reg_10136_pp0_iter3_reg + data_10_V_read11_reg_10105_pp0_iter3_reg);

assign add_ln703_210_fu_1314_p2 = (add_ln703_209_reg_10646 + sub_ln703_68_fu_1133_p2);

assign add_ln703_211_fu_1339_p2 = (sub_ln703_84_fu_1222_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_213_fu_1068_p2 = (sub_ln703_46_fu_858_p2 + data_10_V_read11_reg_10105_pp0_iter3_reg);

assign add_ln703_214_fu_1349_p2 = (add_ln703_213_reg_10653 + data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign add_ln703_215_fu_1353_p2 = (add_ln703_214_fu_1349_p2 + add_ln703_192_reg_10626);

assign add_ln703_216_fu_1358_p2 = (sub_ln703_85_fu_1230_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_217_fu_1393_p2 = (add_ln703_162_reg_10539 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_219_fu_1397_p2 = (add_ln703_209_reg_10646 + add_ln703_217_fu_1393_p2);

assign add_ln703_221_fu_1402_p2 = (add_ln703_209_reg_10646 + sub_ln703_76_fu_1155_p2);

assign add_ln703_222_fu_1626_p2 = (sub_ln703_96_reg_10677 + data_11_V_read12_reg_10075_pp0_iter5_reg);

assign add_ln703_223_fu_1073_p2 = (data_10_V_read11_reg_10105_pp0_iter3_reg + data_11_V_read12_reg_10075_pp0_iter3_reg);

assign add_ln703_224_fu_1437_p2 = (add_ln703_223_reg_10658 + sub_ln703_81_fu_1194_p2);

assign add_ln703_225_fu_1452_p2 = (sub_ln703_102_fu_1344_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_226_fu_1457_p2 = (add_ln703_215_fu_1353_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_227_fu_1472_p2 = (sub_ln703_104_fu_1368_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_228_fu_1477_p2 = (sub_ln703_105_fu_1373_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_229_fu_1654_p2 = (sub_ln703_107_reg_10712 + data_11_V_read12_reg_10075_pp0_iter5_reg);

assign add_ln703_230_fu_1658_p2 = (sub_ln703_108_reg_10717 + data_11_V_read12_reg_10075_pp0_iter5_reg);

assign add_ln703_232_fu_1492_p2 = (add_ln703_223_reg_10658 + sub_ln703_92_reg_10636);

assign add_ln703_233_fu_1501_p2 = (sub_ln703_112_fu_1422_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_234_fu_1671_p2 = (sub_ln703_114_fu_1630_p2 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_235_fu_1676_p2 = (sub_ln703_115_reg_10727 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_236_fu_1511_p2 = (sub_ln703_119_fu_1442_p2 + data_12_V_read13_reg_10045_pp0_iter4_reg);

assign add_ln703_237_fu_1516_p2 = (data_11_V_read12_reg_10075_pp0_iter4_reg + data_12_V_read13_reg_10045_pp0_iter4_reg);

assign add_ln703_238_fu_1520_p2 = (add_ln703_237_fu_1516_p2 + sub_ln703_100_fu_1329_p2);

assign add_ln703_240_fu_1526_p2 = (add_ln703_237_fu_1516_p2 + sub_ln703_101_fu_1334_p2);

assign add_ln703_241_fu_1693_p2 = (sub_ln703_121_fu_1646_p2 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_242_fu_1537_p2 = (sub_ln703_86_fu_1234_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_244_fu_1542_p2 = (add_ln703_237_fu_1516_p2 + add_ln703_242_fu_1537_p2);

assign add_ln703_245_fu_1721_p2 = (sub_ln703_125_reg_10757 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_247_fu_1563_p2 = (add_ln703_237_fu_1516_p2 + sub_ln703_110_fu_1412_p2);

assign add_ln703_248_fu_1569_p2 = (sub_ln703_95_fu_1285_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_250_fu_1574_p2 = (add_ln703_237_fu_1516_p2 + add_ln703_248_fu_1569_p2);

assign add_ln703_251_fu_1753_p2 = (sub_ln703_131_fu_1680_p2 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_252_fu_1077_p2 = (data_12_V_read13_reg_10045_pp0_iter3_reg + data_13_V_read14_reg_10015_pp0_iter3_reg);

assign add_ln703_253_fu_1758_p2 = (add_ln703_252_reg_10665_pp0_iter5_reg + sub_ln703_117_fu_1638_p2);

assign add_ln703_254_fu_1081_p2 = (sub_ln703_42_fu_833_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_256_fu_1585_p2 = (add_ln703_192_reg_10626 + add_ln703_254_reg_10672);

assign add_ln703_259_fu_1589_p2 = (add_ln703_252_reg_10665 + add_ln703_223_reg_10658);

assign add_ln703_260_fu_1593_p2 = (add_ln703_259_fu_1589_p2 + add_ln703_256_fu_1585_p2);

assign add_ln703_262_fu_1604_p2 = (add_ln703_252_reg_10665 + sub_ln703_120_fu_1447_p2);

assign add_ln703_263_fu_1771_p2 = (sub_ln703_133_reg_10782 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_264_fu_1821_p2 = (sub_ln703_145_fu_1734_p2 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_265_fu_1614_p2 = (data_13_V_read14_reg_10015_pp0_iter4_reg + data_14_V_read15_reg_9987_pp0_iter4_reg);

assign add_ln703_266_fu_1854_p2 = (add_ln703_265_reg_10837 + sub_ln703_132_fu_1684_p2);

assign add_ln703_268_fu_1886_p2 = (add_ln703_265_reg_10837 + sub_ln703_134_fu_1689_p2);

assign add_ln703_269_fu_1891_p2 = (sub_ln703_122_reg_10742 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_271_fu_1895_p2 = (add_ln703_265_reg_10837 + add_ln703_269_fu_1891_p2);

assign add_ln703_273_fu_1914_p2 = (add_ln703_265_reg_10837 + sub_ln703_138_fu_1706_p2);

assign add_ln703_274_fu_1924_p2 = (sub_ln703_161_fu_1809_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_276_fu_1934_p2 = (add_ln703_265_reg_10837 + sub_ln703_143_fu_1725_p2);

assign add_ln703_277_fu_1939_p2 = (sub_ln703_163_fu_1817_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_278_fu_1954_p2 = (sub_ln703_165_fu_1830_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_279_fu_1964_p2 = (sub_ln703_116_fu_1634_p2 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_280_fu_1618_p2 = (data_14_V_read15_reg_9987_pp0_iter4_reg + data_15_V_read16_reg_9962_pp0_iter4_reg);

assign add_ln703_281_fu_1969_p2 = (add_ln703_280_reg_10846 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_282_fu_1973_p2 = (add_ln703_281_fu_1969_p2 + add_ln703_279_fu_1964_p2);

assign add_ln703_283_fu_1979_p2 = (sub_ln703_169_fu_1849_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_285_fu_2009_p2 = (add_ln703_280_reg_10846 + sub_ln703_153_fu_1775_p2);

assign add_ln703_287_fu_2019_p2 = (add_ln703_280_reg_10846 + sub_ln703_155_fu_1780_p2);

assign add_ln703_289_fu_2034_p2 = (add_ln703_280_reg_10846 + sub_ln703_158_fu_1794_p2);

assign add_ln703_290_fu_2039_p2 = (sub_ln703_179_fu_1919_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_291_fu_2064_p2 = (sub_ln703_144_fu_1730_p2 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_293_fu_2069_p2 = (add_ln703_280_reg_10846 + add_ln703_291_fu_2064_p2);

assign add_ln703_294_fu_2084_p2 = (sub_ln703_147_fu_1738_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_295_fu_2089_p2 = (data_15_V_read16_reg_9962_pp0_iter5_reg + data_16_V_read17_reg_9935_pp0_iter5_reg);

assign add_ln703_296_fu_2238_p2 = (add_ln703_295_reg_10923 + add_ln703_294_reg_10918);

assign add_ln703_298_fu_2242_p2 = (add_ln703_295_reg_10923 + sub_ln703_166_reg_10863);

assign add_ln703_300_fu_2093_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_167_fu_1839_p2);

assign add_ln703_301_fu_2250_p2 = (sub_ln703_184_reg_10878 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_303_fu_2104_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_171_fu_1864_p2);

assign add_ln703_304_fu_2110_p2 = (sub_ln703_185_fu_1989_p2 + data_16_V_read17_reg_9935_pp0_iter5_reg);

assign add_ln703_305_fu_2254_p2 = (sub_ln703_186_reg_10883 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_307_fu_2125_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_176_fu_1900_p2);

assign add_ln703_309_fu_2136_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_177_fu_1904_p2);

assign add_ln703_310_fu_2147_p2 = (sub_ln703_159_fu_1799_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_312_fu_2270_p2 = (add_ln703_295_reg_10923 + add_ln703_310_reg_10980);

assign add_ln703_314_fu_2167_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_182_fu_1949_p2);

assign add_ln703_315_fu_2300_p2 = (sub_ln703_199_fu_2246_p2 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_316_fu_2178_p2 = (data_16_V_read17_reg_9935_pp0_iter5_reg + data_17_V_read18_reg_9904_pp0_iter5_reg);

assign add_ln703_317_fu_2182_p2 = (add_ln703_316_fu_2178_p2 + sub_ln703_187_fu_1999_p2);

assign add_ln703_318_fu_2323_p2 = (sub_ln703_201_fu_2258_p2 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_319_fu_2328_p2 = (sub_ln703_202_reg_10955 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_320_fu_2336_p2 = (sub_ln703_203_reg_10965 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_321_fu_2353_p2 = (sub_ln703_206_fu_2266_p2 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_323_fu_2188_p2 = (add_ln703_316_fu_2178_p2 + sub_ln703_193_fu_2049_p2);

assign add_ln703_324_fu_2405_p2 = (sub_ln703_217_fu_2305_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_325_fu_2199_p2 = (sub_ln703_170_fu_1859_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_326_fu_1622_p2 = (data_17_V_read18_reg_9904_pp0_iter4_reg + data_18_V_read_8_reg_9874_pp0_iter4_reg);

assign add_ln703_327_fu_2204_p2 = (add_ln703_326_reg_10855 + data_16_V_read17_reg_9935_pp0_iter5_reg);

assign add_ln703_328_fu_2208_p2 = (add_ln703_327_fu_2204_p2 + add_ln703_325_fu_2199_p2);

assign add_ln703_329_fu_2410_p2 = (sub_ln703_218_fu_2310_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_330_fu_2219_p2 = (sub_ln703_175_fu_1881_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_333_fu_2224_p2 = (add_ln703_327_fu_2204_p2 + add_ln703_330_fu_2219_p2);

assign add_ln703_335_fu_2420_p2 = (add_ln703_326_reg_10855_pp0_iter6_reg + sub_ln703_200_reg_10950);

assign add_ln703_336_fu_2449_p2 = (sub_ln703_224_fu_2348_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_337_fu_2459_p2 = (sub_ln703_225_fu_2358_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_339_fu_2464_p2 = (add_ln703_326_reg_10855_pp0_iter6_reg + sub_ln703_208_reg_10985);

assign add_ln703_340_fu_2491_p2 = (sub_ln703_231_fu_2381_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_341_fu_2230_p2 = (data_18_V_read_8_reg_9874_pp0_iter5_reg + data_19_V_read_8_reg_9845_pp0_iter5_reg);

assign add_ln703_342_fu_2520_p2 = (add_ln703_341_reg_11030 + sub_ln703_219_fu_2314_p2);

assign add_ln703_343_fu_2554_p2 = (sub_ln703_241_fu_2439_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_345_fu_2564_p2 = (add_ln703_341_reg_11030 + sub_ln703_223_fu_2344_p2);

assign add_ln703_346_fu_2589_p2 = (sub_ln703_244_fu_2468_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_347_fu_2594_p2 = (sub_ln703_194_reg_10908 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_349_fu_2598_p2 = (add_ln703_341_reg_11030 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_350_fu_2602_p2 = (add_ln703_349_fu_2598_p2 + add_ln703_347_fu_2594_p2);

assign add_ln703_351_fu_2608_p2 = (sub_ln703_245_fu_2472_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_352_fu_2633_p2 = (sub_ln703_253_fu_2515_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_353_fu_2795_p2 = (sub_ln703_254_reg_11076 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_354_fu_2638_p2 = (data_19_V_read_8_reg_9845_pp0_iter6_reg + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_355_fu_2642_p2 = (add_ln703_354_fu_2638_p2 + sub_ln703_237_reg_11020);

assign add_ln703_356_fu_2657_p2 = (sub_ln703_259_fu_2549_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_357_fu_2811_p2 = (sub_ln703_263_reg_11101 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_358_fu_2672_p2 = (sub_ln703_226_fu_2363_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_360_fu_2677_p2 = (add_ln703_354_fu_2638_p2 + add_ln703_358_fu_2672_p2);

assign add_ln703_361_fu_2683_p2 = (sub_ln703_264_fu_2584_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_363_fu_2823_p2 = (add_ln703_354_reg_11131 + sub_ln703_246_reg_11051);

assign add_ln703_364_fu_2831_p2 = (sub_ln703_268_fu_2783_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_365_fu_2841_p2 = (sub_ln703_270_reg_11121 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_366_fu_2871_p2 = (sub_ln703_275_reg_11153 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_367_fu_2903_p2 = (sub_ln703_284_reg_11168 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_368_fu_2723_p2 = (sub_ln703_233_fu_2390_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_369_fu_2234_p2 = (data_21_V_read22_reg_9784_pp0_iter5_reg + data_22_V_read23_reg_9756_pp0_iter5_reg);

assign add_ln703_370_fu_2728_p2 = (add_ln703_369_reg_11037 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_371_fu_2732_p2 = (add_ln703_370_fu_2728_p2 + add_ln703_368_fu_2723_p2);

assign add_ln703_372_fu_2927_p2 = (sub_ln703_289_reg_11173 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_374_fu_2936_p2 = (add_ln703_369_reg_11037_pp0_iter7_reg + sub_ln703_273_fu_2799_p2);

assign add_ln703_375_fu_2738_p2 = (sub_ln703_260_fu_2559_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_377_fu_2956_p2 = (add_ln703_369_reg_11037_pp0_iter7_reg + add_ln703_375_reg_11198);

assign add_ln703_378_fu_2960_p2 = (sub_ln703_293_reg_11178 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_379_fu_2964_p2 = (sub_ln703_295_fu_2880_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_380_fu_2969_p2 = (sub_ln703_296_reg_11183 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_381_fu_2973_p2 = (sub_ln703_297_fu_2884_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_382_fu_2983_p2 = (sub_ln703_299_fu_2894_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_383_fu_3007_p2 = (sub_ln703_250_reg_11061 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_384_fu_2743_p2 = (data_22_V_read23_reg_9756_pp0_iter6_reg + data_23_V_read24_reg_9730_pp0_iter6_reg);

assign add_ln703_385_fu_3011_p2 = (add_ln703_384_reg_11203 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_386_fu_3015_p2 = (add_ln703_385_fu_3011_p2 + add_ln703_383_fu_3007_p2);

assign add_ln703_387_fu_3046_p2 = (sub_ln703_257_reg_11086 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_390_fu_3050_p2 = (add_ln703_385_fu_3011_p2 + add_ln703_387_fu_3046_p2);

assign add_ln703_391_fu_3061_p2 = (sub_ln703_308_fu_2946_p2 + data_23_V_read24_reg_9730_pp0_iter7_reg);

assign add_ln703_392_fu_3081_p2 = (sub_ln703_277_fu_2803_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_394_fu_3086_p2 = (add_ln703_384_reg_11203 + add_ln703_392_fu_3081_p2);

assign add_ln703_395_fu_3116_p2 = (sub_ln703_282_fu_2827_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_397_fu_3121_p2 = (add_ln703_384_reg_11203 + add_ln703_395_fu_3116_p2);

assign add_ln703_398_fu_2747_p2 = (sub_ln703_214_fu_2287_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_400_fu_2752_p2 = (add_ln703_354_fu_2638_p2 + add_ln703_398_fu_2747_p2);

assign add_ln703_402_fu_2758_p2 = (data_23_V_read24_reg_9730_pp0_iter6_reg + data_24_V_read25_reg_9704_pp0_iter6_reg);

assign add_ln703_403_fu_3131_p2 = (add_ln703_402_reg_11215 + add_ln703_369_reg_11037_pp0_iter7_reg);

assign add_ln703_404_fu_3135_p2 = (add_ln703_403_fu_3131_p2 + add_ln703_400_reg_11210);

assign add_ln703_406_fu_3145_p2 = (add_ln703_354_reg_11131 + sub_ln703_234_reg_11046);

assign add_ln703_410_fu_3149_p2 = (add_ln703_403_fu_3131_p2 + add_ln703_406_fu_3145_p2);

assign add_ln703_411_fu_3380_p2 = (sub_ln703_315_reg_11267 + data_24_V_read25_reg_9704_pp0_iter8_reg);

assign add_ln703_413_fu_3160_p2 = (add_ln703_402_reg_11215 + sub_ln703_305_fu_2922_p2);

assign add_ln703_414_fu_3165_p2 = (sub_ln703_288_fu_2854_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_416_fu_3170_p2 = (add_ln703_402_reg_11215 + add_ln703_414_fu_3165_p2);

assign add_ln703_417_fu_3185_p2 = (sub_ln703_321_fu_3066_p2 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_418_fu_3210_p2 = (sub_ln703_325_fu_3096_p2 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_419_fu_3225_p2 = (sub_ln703_301_reg_11188 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_421_fu_3229_p2 = (add_ln703_402_reg_11215 + add_ln703_419_fu_3225_p2);

assign add_ln703_422_fu_3239_p2 = (sub_ln703_331_fu_3140_p2 + data_25_V_read26_reg_9677_pp0_iter7_reg);

assign add_ln703_423_fu_3249_p2 = (sub_ln703_287_fu_2849_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_424_fu_2762_p2 = (data_24_V_read25_reg_9704_pp0_iter6_reg + data_25_V_read26_reg_9677_pp0_iter6_reg);

assign add_ln703_425_fu_3254_p2 = (add_ln703_424_reg_11225 + data_23_V_read24_reg_9730_pp0_iter7_reg);

assign add_ln703_426_fu_3258_p2 = (add_ln703_425_fu_3254_p2 + add_ln703_423_fu_3249_p2);

assign add_ln703_428_fu_3264_p2 = (add_ln703_424_reg_11225 + sub_ln703_317_fu_3031_p2);

assign add_ln703_429_fu_3418_p2 = (sub_ln703_335_fu_3384_p2 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_430_fu_3423_p2 = (sub_ln703_336_reg_11307 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_431_fu_3274_p2 = (sub_ln703_338_fu_3195_p2 + data_25_V_read26_reg_9677_pp0_iter7_reg);

assign add_ln703_432_fu_3279_p2 = (sub_ln703_294_fu_2875_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_435_fu_3284_p2 = (add_ln703_425_fu_3254_p2 + add_ln703_432_fu_3279_p2);

assign add_ln703_436_fu_3439_p2 = (sub_ln703_342_reg_11327 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_437_fu_3443_p2 = (sub_ln703_346_fu_3396_p2 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_438_fu_3310_p2 = (sub_ln703_320_fu_3056_p2 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_439_fu_2766_p2 = (data_25_V_read26_reg_9677_pp0_iter6_reg + data_26_V_read27_reg_9652_pp0_iter6_reg);

assign add_ln703_440_fu_3466_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + add_ln703_438_reg_11382);

assign add_ln703_441_fu_3480_p2 = (sub_ln703_353_reg_11352 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_442_fu_3502_p2 = (sub_ln703_356_reg_11367 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_444_fu_3506_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + sub_ln703_341_fu_3388_p2);

assign add_ln703_445_fu_3315_p2 = (sub_ln703_310_fu_2978_p2 + data_23_V_read24_reg_9730_pp0_iter7_reg);

assign add_ln703_447_fu_3320_p2 = (add_ln703_439_reg_11233 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_448_fu_3511_p2 = (add_ln703_447_reg_11392 + add_ln703_445_reg_11387);

assign add_ln703_450_fu_3520_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + sub_ln703_344_reg_11332);

assign add_ln703_451_fu_3329_p2 = (data_26_V_read27_reg_9652_pp0_iter7_reg + data_27_V_read28_reg_9625_pp0_iter7_reg);

assign add_ln703_452_fu_3524_p2 = (add_ln703_451_reg_11402 + sub_ln703_345_reg_11337);

assign add_ln703_453_fu_3528_p2 = (sub_ln703_358_reg_11372 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_455_fu_3537_p2 = (add_ln703_451_reg_11402 + sub_ln703_348_fu_3405_p2);

assign add_ln703_456_fu_3542_p2 = (sub_ln703_359_fu_3448_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_458_fu_3552_p2 = (add_ln703_451_reg_11402 + sub_ln703_351_fu_3414_p2);

assign add_ln703_459_fu_3557_p2 = (sub_ln703_334_reg_11302 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_461_fu_3561_p2 = (add_ln703_451_reg_11402 + add_ln703_459_fu_3557_p2);

assign add_ln703_462_fu_3571_p2 = (sub_ln703_364_fu_3470_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_463_fu_3581_p2 = (sub_ln703_366_fu_3484_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_464_fu_3586_p2 = (sub_ln703_367_fu_3488_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_465_fu_3630_p2 = (sub_ln703_330_fu_3372_p2 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_466_fu_3333_p2 = (data_27_V_read28_reg_9625_pp0_iter7_reg + data_28_V_read_8_reg_9598_pp0_iter7_reg);

assign add_ln703_467_fu_3635_p2 = (add_ln703_466_reg_11410 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_468_fu_3639_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_465_fu_3630_p2);

assign add_ln703_469_fu_3655_p2 = (sub_ln703_372_fu_3532_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_471_fu_3337_p2 = (add_ln703_424_reg_11225 + sub_ln703_319_fu_3041_p2);

assign add_ln703_474_fu_3680_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_471_reg_11418);

assign add_ln703_476_fu_3685_p2 = (add_ln703_466_reg_11410 + sub_ln703_363_fu_3461_p2);

assign add_ln703_477_fu_3715_p2 = (sub_ln703_378_fu_3601_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_478_fu_3730_p2 = (sub_ln703_381_fu_3616_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_479_fu_3735_p2 = (sub_ln703_343_fu_3392_p2 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_482_fu_3740_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_479_fu_3735_p2);

assign add_ln703_484_fu_3342_p2 = (add_ln703_424_reg_11225 + sub_ln703_329_fu_3126_p2);

assign add_ln703_487_fu_3756_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_484_reg_11423);

assign add_ln703_488_fu_3766_p2 = (sub_ln703_385_fu_3650_p2 + data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign add_ln703_489_fu_3771_p2 = (sub_ln703_361_fu_3457_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_490_fu_3347_p2 = (data_28_V_read_8_reg_9598_pp0_iter7_reg + data_29_V_read_8_reg_9573_pp0_iter7_reg);

assign add_ln703_491_fu_3776_p2 = (add_ln703_490_reg_11428 + add_ln703_489_fu_3771_p2);

assign add_ln703_493_fu_3796_p2 = (add_ln703_490_reg_11428 + sub_ln703_374_fu_3566_p2);

assign add_ln703_494_fu_3801_p2 = (sub_ln703_365_fu_3475_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_496_fu_3806_p2 = (add_ln703_490_reg_11428 + add_ln703_494_fu_3801_p2);

assign add_ln703_497_fu_3811_p2 = (sub_ln703_391_fu_3695_p2 + data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign add_ln703_498_fu_3351_p2 = (sub_ln703_278_fu_2807_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_500_fu_3821_p2 = (add_ln703_402_reg_11215_pp0_iter8_reg + data_22_V_read23_reg_9756_pp0_iter8_reg);

assign add_ln703_501_fu_3825_p2 = (add_ln703_500_fu_3821_p2 + add_ln703_498_reg_11436);

assign add_ln703_504_fu_3830_p2 = (add_ln703_490_reg_11428 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_505_fu_3834_p2 = (add_ln703_504_fu_3830_p2 + add_ln703_439_reg_11233_pp0_iter8_reg);

assign add_ln703_506_fu_3839_p2 = (add_ln703_505_fu_3834_p2 + add_ln703_501_fu_3825_p2);

assign add_ln703_507_fu_3356_p2 = (data_29_V_read_8_reg_9573_pp0_iter7_reg + data_30_V_read31_reg_9549_pp0_iter7_reg);

assign add_ln703_508_fu_4006_p2 = (add_ln703_507_reg_11441_pp0_iter9_reg + sub_ln703_386_reg_11484);

assign add_ln703_509_fu_3870_p2 = (sub_ln703_362_reg_11377 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_511_fu_3874_p2 = (add_ln703_507_reg_11441 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_512_fu_3878_p2 = (add_ln703_511_fu_3874_p2 + add_ln703_509_fu_3870_p2);

assign add_ln703_513_fu_4035_p2 = (sub_ln703_407_fu_3985_p2 + data_30_V_read31_reg_9549_pp0_iter9_reg);

assign add_ln703_515_fu_3889_p2 = (add_ln703_507_reg_11441 + sub_ln703_396_fu_3725_p2);

assign add_ln703_517_fu_3894_p2 = (add_ln703_507_reg_11441 + sub_ln703_397_fu_3746_p2);

assign add_ln703_519_fu_3899_p2 = (add_ln703_507_reg_11441 + sub_ln703_398_fu_3751_p2);

assign add_ln703_520_fu_4058_p2 = (sub_ln703_412_reg_11574 + data_30_V_read31_reg_9549_pp0_iter9_reg);

assign add_ln703_521_fu_4062_p2 = (sub_ln703_413_fu_3997_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_522_fu_4067_p2 = (sub_ln703_414_reg_11579 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_523_fu_2770_p2 = (sub_ln703_183_reg_10868 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_525_fu_2774_p2 = (add_ln703_326_reg_10855_pp0_iter6_reg + add_ln703_523_fu_2770_p2);

assign add_ln703_528_fu_3360_p2 = (add_ln703_369_reg_11037_pp0_iter7_reg + add_ln703_354_reg_11131);

assign add_ln703_529_fu_4071_p2 = (add_ln703_528_reg_11452_pp0_iter9_reg + add_ln703_525_reg_11243_pp0_iter9_reg);

assign add_ln703_532_fu_3904_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + add_ln703_402_reg_11215_pp0_iter8_reg);

assign add_ln703_534_fu_2779_p2 = (data_30_V_read31_reg_9549_pp0_iter6_reg + data_31_V_read32_reg_9521_pp0_iter6_reg);

assign add_ln703_535_fu_3364_p2 = (add_ln703_534_reg_11248 + data_29_V_read_8_reg_9573_pp0_iter7_reg);

assign add_ln703_536_fu_3908_p2 = (add_ln703_535_reg_11457 + add_ln703_466_reg_11410);

assign add_ln703_537_fu_3912_p2 = (add_ln703_536_fu_3908_p2 + add_ln703_532_fu_3904_p2);

assign add_ln703_538_fu_4075_p2 = (add_ln703_537_reg_11609 + add_ln703_529_fu_4071_p2);

assign add_ln703_539_fu_4085_p2 = (sub_ln703_387_reg_11489 + data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign add_ln703_541_fu_4089_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + add_ln703_539_fu_4085_p2);

assign add_ln703_542_fu_3918_p2 = (sub_ln703_373_fu_3547_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_545_fu_3923_p2 = (add_ln703_535_reg_11457 + add_ln703_542_fu_3918_p2);

assign add_ln703_546_fu_4094_p2 = (sub_ln703_416_reg_11584 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_548_fu_4098_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + sub_ln703_401_reg_11529);

assign add_ln703_550_fu_4111_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + sub_ln703_403_reg_11539);

assign add_ln703_551_fu_4115_p2 = (sub_ln703_418_fu_4014_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_552_fu_4139_p2 = (sub_ln703_423_fu_4031_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_553_fu_3928_p2 = (sub_ln703_376_fu_3591_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_556_fu_3933_p2 = (add_ln703_535_reg_11457 + add_ln703_553_fu_3928_p2);

assign add_ln703_557_fu_4158_p2 = (sub_ln703_426_fu_4049_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_558_fu_4216_p2 = (sub_ln703_429_fu_4102_p2 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_559_fu_4241_p2 = (sub_ln703_432_fu_4124_p2 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_560_fu_3943_p2 = (data_31_V_read32_reg_9521_pp0_iter8_reg + data_32_V_read_3_reg_9492_pp0_iter8_reg);

assign add_ln703_561_fu_4260_p2 = (add_ln703_560_reg_11629 + sub_ln703_425_fu_4044_p2);

assign add_ln703_562_fu_4275_p2 = (sub_ln703_439_fu_4168_p2 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_563_fu_4280_p2 = (sub_ln703_440_reg_11624 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_564_fu_3947_p2 = (sub_ln703_347_fu_3400_p2 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_566_fu_3952_p2 = (add_ln703_466_reg_11410 + add_ln703_564_fu_3947_p2);

assign add_ln703_568_fu_3368_p2 = (data_32_V_read_3_reg_9492_pp0_iter7_reg + data_33_V_read_3_reg_9463_pp0_iter7_reg);

assign add_ln703_569_fu_3957_p2 = (add_ln703_568_reg_11464 + data_31_V_read32_reg_9521_pp0_iter8_reg);

assign add_ln703_570_fu_4294_p2 = (add_ln703_569_reg_11640 + add_ln703_507_reg_11441_pp0_iter9_reg);

assign add_ln703_571_fu_4298_p2 = (add_ln703_570_fu_4294_p2 + add_ln703_566_reg_11635);

assign add_ln703_572_fu_4308_p2 = (sub_ln703_446_fu_4197_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_573_fu_4323_p2 = (sub_ln703_450_fu_4221_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_574_fu_4566_p2 = (sub_ln703_453_reg_11683 + data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign add_ln703_576_fu_4338_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_433_fu_4129_p2);

assign add_ln703_577_fu_4343_p2 = (sub_ln703_406_fu_3981_p2 + data_30_V_read31_reg_9549_pp0_iter9_reg);

assign add_ln703_580_fu_4348_p2 = (add_ln703_569_reg_11640 + add_ln703_577_fu_4343_p2);

assign add_ln703_581_fu_4358_p2 = (sub_ln703_455_fu_4251_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_583_fu_4363_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_435_fu_4144_p2);

assign add_ln703_585_fu_4383_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_438_fu_4163_p2);

assign add_ln703_586_fu_4398_p2 = (sub_ln703_460_fu_4289_p2 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_587_fu_4403_p2 = (sub_ln703_415_fu_4001_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_588_fu_3961_p2 = (data_33_V_read_3_reg_9463_pp0_iter8_reg + data_34_V_read_3_reg_9434_pp0_iter8_reg);

assign add_ln703_589_fu_4408_p2 = (add_ln703_588_reg_11646 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_590_fu_4412_p2 = (add_ln703_589_fu_4408_p2 + add_ln703_587_fu_4403_p2);

assign add_ln703_591_fu_4423_p2 = (sub_ln703_464_fu_4318_p2 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_592_fu_4428_p2 = (sub_ln703_465_fu_4328_p2 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_594_fu_4433_p2 = (add_ln703_507_reg_11441_pp0_iter9_reg + sub_ln703_390_reg_11499);

assign add_ln703_597_fu_4437_p2 = (add_ln703_588_reg_11646 + add_ln703_560_reg_11629);

assign add_ln703_598_fu_4441_p2 = (add_ln703_597_fu_4437_p2 + add_ln703_594_fu_4433_p2);

assign add_ln703_599_fu_4477_p2 = (sub_ln703_442_fu_4177_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_600_fu_3965_p2 = (data_34_V_read_3_reg_9434_pp0_iter8_reg + data_35_V_read_3_reg_9410_pp0_iter8_reg);

assign add_ln703_601_fu_4620_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + add_ln703_599_reg_11798);

assign add_ln703_602_fu_4482_p2 = (sub_ln703_384_reg_11474 + data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign add_ln703_604_fu_4486_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + add_ln703_602_fu_4482_p2);

assign add_ln703_607_fu_4491_p2 = (add_ln703_600_reg_11652 + add_ln703_568_reg_11464_pp0_iter9_reg);

assign add_ln703_608_fu_4495_p2 = (add_ln703_607_fu_4491_p2 + add_ln703_604_fu_4486_p2);

assign add_ln703_609_fu_4501_p2 = (sub_ln703_444_fu_4187_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_611_fu_4628_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + add_ln703_609_reg_11803);

assign add_ln703_612_fu_4640_p2 = (sub_ln703_477_fu_4578_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_613_fu_4645_p2 = (sub_ln703_478_fu_4582_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_614_fu_4506_p2 = (sub_ln703_449_fu_4211_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_616_fu_4511_p2 = (add_ln703_600_reg_11652 + add_ln703_614_fu_4506_p2);

assign add_ln703_617_fu_4677_p2 = (sub_ln703_484_fu_4599_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_618_fu_4687_p2 = (sub_ln703_486_fu_4607_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_619_fu_4692_p2 = (sub_ln703_488_reg_11783 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_620_fu_4696_p2 = (sub_ln703_491_reg_11793 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_621_fu_3969_p2 = (data_35_V_read_3_reg_9410_pp0_iter8_reg + data_36_V_read_3_reg_9383_pp0_iter8_reg);

assign add_ln703_622_fu_4720_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_476_fu_4574_p2);

assign add_ln703_623_fu_4739_p2 = (sub_ln703_496_fu_4650_p2 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_624_fu_4754_p2 = (sub_ln703_466_fu_4562_p2 + data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign add_ln703_626_fu_4759_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + add_ln703_624_fu_4754_p2);

assign add_ln703_627_fu_4769_p2 = (sub_ln703_501_fu_4672_p2 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_629_fu_4774_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_482_reg_11773);

assign add_ln703_631_fu_4526_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_434_fu_4134_p2);

assign add_ln703_633_fu_4531_p2 = (add_ln703_621_reg_11662 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_634_fu_4535_p2 = (add_ln703_633_fu_4531_p2 + add_ln703_631_fu_4526_p2);

assign add_ln703_636_fu_4793_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_487_fu_4611_p2);

assign add_ln703_638_fu_4803_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_489_fu_4615_p2);

assign add_ln703_639_fu_4541_p2 = (sub_ln703_459_fu_4284_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_642_fu_4817_p2 = (add_ln703_633_reg_11823 + add_ln703_639_reg_11833);

assign add_ln703_643_fu_4821_p2 = (sub_ln703_504_fu_4700_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_644_fu_4826_p2 = (sub_ln703_505_reg_11818 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_645_fu_4835_p2 = (sub_ln703_507_fu_4710_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_646_fu_4546_p2 = (data_36_V_read_3_reg_9383_pp0_iter9_reg + data_37_V_read_3_reg_9353_pp0_iter9_reg);

assign add_ln703_647_fu_4870_p2 = (add_ln703_646_reg_11838 + sub_ln703_499_fu_4663_p2);

assign add_ln703_648_fu_4899_p2 = (sub_ln703_516_fu_4783_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_649_fu_4914_p2 = (sub_ln703_518_fu_4798_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_650_fu_4550_p2 = (data_37_V_read_3_reg_9353_pp0_iter9_reg + data_38_V_read_3_reg_9328_pp0_iter9_reg);

assign add_ln703_651_fu_4959_p2 = (add_ln703_650_reg_11844 + sub_ln703_510_fu_4730_p2);

assign add_ln703_653_fu_4964_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + sub_ln703_463_fu_4558_p2);

assign add_ln703_655_fu_4969_p2 = (add_ln703_650_reg_11844 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_656_fu_4973_p2 = (add_ln703_655_fu_4969_p2 + add_ln703_653_fu_4964_p2);

assign add_ln703_658_fu_4989_p2 = (add_ln703_650_reg_11844 + sub_ln703_513_fu_4749_p2);

assign add_ln703_659_fu_5150_p2 = (sub_ln703_529_reg_11879 + data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign add_ln703_660_fu_4994_p2 = (sub_ln703_531_fu_4890_p2 + data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign add_ln703_661_fu_4999_p2 = (sub_ln703_534_fu_4909_p2 + data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign add_ln703_662_fu_5166_p2 = (sub_ln703_535_reg_11899 + data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign add_ln703_663_fu_5009_p2 = (sub_ln703_490_reg_11788 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_666_fu_5013_p2 = (add_ln703_655_fu_4969_p2 + add_ln703_663_fu_5009_p2);

assign add_ln703_667_fu_4554_p2 = (data_38_V_read_3_reg_9328_pp0_iter9_reg + data_39_V_read_3_reg_9301_pp0_iter9_reg);

assign add_ln703_668_fu_5019_p2 = (add_ln703_667_reg_11853 + sub_ln703_521_fu_4830_p2);

assign add_ln703_669_fu_5186_p2 = (sub_ln703_544_reg_11934 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_671_fu_5039_p2 = (add_ln703_667_reg_11853 + sub_ln703_530_fu_4885_p2);

assign add_ln703_673_fu_5044_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_483_reg_11778);

assign add_ln703_675_fu_5048_p2 = (add_ln703_667_reg_11853 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_676_fu_5052_p2 = (add_ln703_675_fu_5048_p2 + add_ln703_673_fu_5044_p2);

assign add_ln703_678_fu_5058_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + sub_ln703_469_reg_11733);

assign add_ln703_681_fu_5062_p2 = (add_ln703_667_reg_11853 + add_ln703_646_reg_11838);

assign add_ln703_682_fu_5066_p2 = (add_ln703_681_fu_5062_p2 + add_ln703_678_fu_5058_p2);

assign add_ln703_683_fu_5072_p2 = (sub_ln703_519_fu_4808_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_685_fu_5077_p2 = (add_ln703_667_reg_11853 + add_ln703_683_fu_5072_p2);

assign add_ln703_687_fu_5082_p2 = (add_ln703_667_reg_11853 + sub_ln703_536_fu_4924_p2);

assign add_ln703_689_fu_5087_p2 = (add_ln703_667_reg_11853 + sub_ln703_537_fu_4929_p2);

assign add_ln703_690_fu_5240_p2 = (sub_ln703_553_fu_5174_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_691_fu_5092_p2 = (data_39_V_read_3_reg_9301_pp0_iter10_reg + data_40_V_read41_reg_9272_pp0_iter10_reg);

assign add_ln703_692_fu_5245_p2 = (add_ln703_691_reg_11994 + sub_ln703_541_reg_11919);

assign add_ln703_693_fu_5249_p2 = (sub_ln703_554_fu_5178_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_694_fu_5254_p2 = (sub_ln703_555_fu_5182_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_695_fu_5259_p2 = (sub_ln703_556_reg_11964 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_696_fu_5272_p2 = (sub_ln703_558_reg_11974 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_697_fu_5096_p2 = (sub_ln703_528_fu_4875_p2 + data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign add_ln703_699_fu_5281_p2 = (add_ln703_691_reg_11994 + add_ln703_697_reg_12002);

assign add_ln703_700_fu_5285_p2 = (sub_ln703_561_fu_5200_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_701_fu_5313_p2 = (sub_ln703_566_fu_5223_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_702_fu_5332_p2 = (sub_ln703_538_reg_11904 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_703_fu_5116_p2 = (data_40_V_read41_reg_9272_pp0_iter10_reg + data_41_V_read42_reg_9242_pp0_iter10_reg);

assign add_ln703_704_fu_5336_p2 = (add_ln703_703_reg_12022 + add_ln703_702_fu_5332_p2);

assign add_ln703_706_fu_5120_p2 = (add_ln703_650_reg_11844 + sub_ln703_509_fu_4725_p2);

assign add_ln703_708_fu_5361_p2 = (add_ln703_703_reg_12022 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_709_fu_5365_p2 = (add_ln703_708_fu_5361_p2 + add_ln703_706_reg_12031);

assign add_ln703_710_fu_5390_p2 = (sub_ln703_545_fu_5138_p2 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_712_fu_5395_p2 = (add_ln703_703_reg_12022 + add_ln703_710_fu_5390_p2);

assign add_ln703_714_fu_5405_p2 = (add_ln703_703_reg_12022 + sub_ln703_559_fu_5190_p2);

assign add_ln703_715_fu_5425_p2 = (sub_ln703_573_reg_12007 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_716_fu_5429_p2 = (sub_ln703_574_fu_5290_p2 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_718_fu_5434_p2 = (add_ln703_703_reg_12022 + sub_ln703_563_fu_5209_p2);

assign add_ln703_719_fu_5439_p2 = (sub_ln703_576_fu_5299_p2 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_720_fu_5469_p2 = (sub_ln703_582_reg_12012 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_721_fu_5692_p2 = (sub_ln703_586_reg_12061 + data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign add_ln703_722_fu_5125_p2 = (sub_ln703_495_fu_4636_p2 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_724_fu_5477_p2 = (add_ln703_650_reg_11844_pp0_iter11_reg + add_ln703_722_reg_12036);

assign add_ln703_726_fu_5130_p2 = (data_41_V_read42_reg_9242_pp0_iter10_reg + data_42_V_read_3_reg_9212_pp0_iter10_reg);

assign add_ln703_727_fu_5481_p2 = (add_ln703_726_reg_12041 + add_ln703_691_reg_11994);

assign add_ln703_728_fu_5485_p2 = (add_ln703_727_fu_5481_p2 + add_ln703_724_fu_5477_p2);

assign add_ln703_729_fu_5700_p2 = (sub_ln703_593_reg_12071 + data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign add_ln703_730_fu_5541_p2 = (sub_ln703_596_fu_5444_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_732_fu_5546_p2 = (add_ln703_726_reg_12041 + sub_ln703_578_fu_5308_p2);

assign add_ln703_733_fu_5551_p2 = (sub_ln703_597_fu_5449_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_734_fu_5556_p2 = (sub_ln703_599_fu_5459_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_735_fu_5571_p2 = (sub_ln703_601_fu_5473_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_736_fu_5576_p2 = (sub_ln703_552_fu_5170_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_737_fu_5134_p2 = (data_42_V_read_3_reg_9212_pp0_iter10_reg + data_43_V_read_3_reg_9184_pp0_iter10_reg);

assign add_ln703_738_fu_5581_p2 = (add_ln703_737_reg_12047 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_739_fu_5585_p2 = (add_ln703_738_fu_5581_p2 + add_ln703_736_fu_5576_p2);

assign add_ln703_741_fu_5591_p2 = (add_ln703_737_reg_12047 + sub_ln703_584_fu_5341_p2);

assign add_ln703_742_fu_5738_p2 = (sub_ln703_605_reg_12111 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_744_fu_5601_p2 = (add_ln703_737_reg_12047 + sub_ln703_592_fu_5400_p2);

assign add_ln703_745_fu_5606_p2 = (sub_ln703_575_fu_5295_p2 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_747_fu_5611_p2 = (add_ln703_737_reg_12047 + add_ln703_745_fu_5606_p2);

assign add_ln703_748_fu_5759_p2 = (sub_ln703_614_reg_12141 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_750_fu_5616_p2 = (add_ln703_691_reg_11994 + sub_ln703_549_fu_5158_p2);

assign add_ln703_753_fu_5621_p2 = (add_ln703_738_fu_5581_p2 + add_ln703_750_fu_5616_p2);

assign add_ln703_754_fu_5776_p2 = (sub_ln703_618_reg_12156 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_755_fu_5652_p2 = (data_43_V_read_3_reg_9184_pp0_iter11_reg + data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign add_ln703_756_fu_5809_p2 = (add_ln703_755_reg_12196 + sub_ln703_606_fu_5696_p2);

assign add_ln703_757_fu_5814_p2 = (sub_ln703_624_reg_12166 + data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign add_ln703_759_fu_5818_p2 = (add_ln703_755_reg_12196 + sub_ln703_608_reg_12116);

assign add_ln703_761_fu_5837_p2 = (add_ln703_755_reg_12196 + sub_ln703_611_fu_5704_p2);

assign add_ln703_763_fu_5842_p2 = (add_ln703_755_reg_12196 + sub_ln703_612_reg_12131);

assign add_ln703_764_fu_5861_p2 = (sub_ln703_630_reg_12171 + data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign add_ln703_765_fu_5671_p2 = (data_44_V_read_3_reg_9154_pp0_iter11_reg + data_45_V_read_3_reg_9125_pp0_iter11_reg);

assign add_ln703_766_fu_5893_p2 = (add_ln703_765_reg_12219 + sub_ln703_621_fu_5726_p2);

assign add_ln703_767_fu_5942_p2 = (sub_ln703_595_reg_12081 + data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign add_ln703_769_fu_5946_p2 = (add_ln703_765_reg_12219 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_770_fu_5950_p2 = (add_ln703_769_fu_5946_p2 + add_ln703_767_fu_5942_p2);

assign add_ln703_771_fu_5961_p2 = (sub_ln703_647_fu_5846_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_772_fu_5966_p2 = (sub_ln703_649_fu_5851_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_774_fu_5985_p2 = (add_ln703_765_reg_12219 + sub_ln703_631_reg_12176);

assign add_ln703_775_fu_5994_p2 = (sub_ln703_616_fu_5712_p2 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_777_fu_5999_p2 = (add_ln703_765_reg_12219 + add_ln703_775_fu_5994_p2);

assign add_ln703_778_fu_5675_p2 = (data_45_V_read_3_reg_9125_pp0_iter11_reg + data_46_V_read_3_reg_9094_pp0_iter11_reg);

assign add_ln703_779_fu_6024_p2 = (add_ln703_778_reg_12227 + sub_ln703_636_fu_5784_p2);

assign add_ln703_781_fu_6029_p2 = (add_ln703_778_reg_12227 + sub_ln703_637_reg_12186);

assign add_ln703_783_fu_5679_p2 = (add_ln703_737_reg_12047 + sub_ln703_585_fu_5346_p2);

assign add_ln703_785_fu_6038_p2 = (add_ln703_778_reg_12227 + data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign add_ln703_786_fu_6042_p2 = (add_ln703_785_fu_6038_p2 + add_ln703_783_reg_12236);

assign add_ln703_788_fu_6082_p2 = (add_ln703_778_reg_12227 + sub_ln703_648_reg_12209);

assign add_ln703_789_fu_6250_p2 = (sub_ln703_669_reg_12268 + data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign add_ln703_790_fu_6121_p2 = (sub_ln703_673_fu_6009_p2 + data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign add_ln703_791_fu_6131_p2 = (sub_ln703_675_fu_6019_p2 + data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign add_ln703_792_fu_6146_p2 = (sub_ln703_677_fu_6047_p2 + data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign add_ln703_793_fu_6258_p2 = (sub_ln703_678_reg_12283 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_794_fu_6151_p2 = (sub_ln703_641_fu_5799_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_795_fu_6156_p2 = (data_46_V_read_3_reg_9094_pp0_iter12_reg + data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign add_ln703_796_fu_6160_p2 = (add_ln703_795_fu_6156_p2 + add_ln703_794_fu_6151_p2);

assign add_ln703_797_fu_6262_p2 = (sub_ln703_681_fu_6238_p2 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_798_fu_6166_p2 = (add_ln703_795_fu_6156_p2 + sub_ln703_663_fu_5923_p2);

assign add_ln703_799_fu_6276_p2 = (sub_ln703_685_fu_6246_p2 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_800_fu_6315_p2 = (sub_ln703_697_reg_12358 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_801_fu_6187_p2 = (sub_ln703_639_fu_5789_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_802_fu_6192_p2 = (data_47_V_read_3_reg_9066_pp0_iter12_reg + data_48_V_read_3_reg_9040_pp0_iter12_reg);

assign add_ln703_803_fu_6319_p2 = (add_ln703_802_reg_12398 + data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign add_ln703_804_fu_6323_p2 = (add_ln703_803_fu_6319_p2 + add_ln703_801_reg_12393);

assign add_ln703_805_fu_6341_p2 = (add_ln703_802_reg_12398 + sub_ln703_680_reg_12293);

assign add_ln703_806_fu_6359_p2 = (sub_ln703_699_fu_6271_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_807_fu_6369_p2 = (sub_ln703_667_reg_12263 + data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign add_ln703_808_fu_6373_p2 = (add_ln703_802_reg_12398 + add_ln703_807_fu_6369_p2);

assign add_ln703_809_fu_6378_p2 = (add_ln703_802_reg_12398 + sub_ln703_686_reg_12308);

assign add_ln703_810_fu_6396_p2 = (sub_ln703_703_fu_6289_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_811_fu_6401_p2 = (sub_ln703_704_reg_12383 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_812_fu_6405_p2 = (add_ln703_802_reg_12398 + sub_ln703_690_reg_12323);

assign add_ln703_813_fu_6409_p2 = (add_ln703_802_reg_12398 + sub_ln703_692_reg_12333);

assign add_ln703_814_fu_6417_p2 = (sub_ln703_708_fu_6302_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_815_fu_6196_p2 = (sub_ln703_661_fu_5913_p2 + data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign add_ln703_816_fu_5684_p2 = (data_48_V_read_3_reg_9040_pp0_iter11_reg + data_49_V_read_3_reg_9012_pp0_iter11_reg);

assign add_ln703_817_fu_6201_p2 = (add_ln703_816_reg_12241 + data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign add_ln703_818_fu_6205_p2 = (add_ln703_817_fu_6201_p2 + add_ln703_815_fu_6196_p2);

assign add_ln703_819_fu_6447_p2 = (sub_ln703_714_fu_6345_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_820_fu_6211_p2 = (add_ln703_778_reg_12227 + sub_ln703_645_fu_5827_p2);

assign add_ln703_821_fu_6216_p2 = (add_ln703_817_fu_6201_p2 + add_ln703_820_fu_6211_p2);

assign add_ln703_822_fu_6482_p2 = (sub_ln703_720_fu_6391_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_823_fu_6512_p2 = (sub_ln703_694_reg_12343 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_824_fu_6516_p2 = (add_ln703_816_reg_12241_pp0_iter13_reg + add_ln703_823_fu_6512_p2);

assign add_ln703_825_fu_6526_p2 = (sub_ln703_722_fu_6422_p2 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_826_fu_6222_p2 = (data_49_V_read_3_reg_9012_pp0_iter12_reg + data_50_V_read51_reg_8984_pp0_iter12_reg);

assign add_ln703_827_fu_6531_p2 = (add_ln703_826_reg_12419 + sub_ln703_710_fu_6311_p2);

assign add_ln703_828_fu_6536_p2 = (add_ln703_826_reg_12419 + sub_ln703_712_fu_6332_p2);

assign add_ln703_829_fu_6546_p2 = (sub_ln703_679_reg_12288 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_830_fu_6550_p2 = (add_ln703_826_reg_12419 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_831_fu_6554_p2 = (add_ln703_830_fu_6550_p2 + add_ln703_829_fu_6546_p2);

assign add_ln703_832_fu_6569_p2 = (sub_ln703_684_reg_12303 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_833_fu_6573_p2 = (add_ln703_830_fu_6550_p2 + add_ln703_832_fu_6569_p2);

assign add_ln703_834_fu_6594_p2 = (sub_ln703_732_fu_6477_p2 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_835_fu_6815_p2 = (sub_ln703_736_reg_12475 + data_50_V_read51_reg_8984_pp0_iter14_reg);

assign add_ln703_836_fu_6226_p2 = (data_50_V_read51_reg_8984_pp0_iter12_reg + data_51_V_read52_reg_8956_pp0_iter12_reg);

assign add_ln703_837_fu_6624_p2 = (add_ln703_836_reg_12428 + sub_ln703_723_fu_6427_p2);

assign add_ln703_838_fu_6634_p2 = (sub_ln703_739_fu_6541_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_839_fu_6836_p2 = (sub_ln703_743_fu_6803_p2 + data_51_V_read52_reg_8956_pp0_iter14_reg);

assign add_ln703_840_fu_6649_p2 = (sub_ln703_747_fu_6584_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_841_fu_6664_p2 = (sub_ln703_752_fu_6609_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_842_fu_6669_p2 = (sub_ln703_705_fu_6294_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_843_fu_6674_p2 = (add_ln703_836_reg_12428 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_844_fu_6678_p2 = (add_ln703_843_fu_6674_p2 + add_ln703_842_fu_6669_p2);

assign add_ln703_845_fu_6689_p2 = (sub_ln703_754_fu_6619_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_846_fu_6863_p2 = (sub_ln703_755_fu_6819_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_847_fu_6868_p2 = (sub_ln703_756_fu_6823_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_848_fu_6694_p2 = (add_ln703_802_reg_12398 + sub_ln703_676_reg_12278);

assign add_ln703_849_fu_6230_p2 = (data_51_V_read52_reg_8956_pp0_iter12_reg + data_52_V_read_3_reg_8928_pp0_iter12_reg);

assign add_ln703_850_fu_6698_p2 = (add_ln703_849_reg_12434 + add_ln703_826_reg_12419);

assign add_ln703_851_fu_6702_p2 = (add_ln703_850_fu_6698_p2 + add_ln703_848_fu_6694_p2);

assign add_ln703_852_fu_6713_p2 = (sub_ln703_711_fu_6328_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_853_fu_6718_p2 = (add_ln703_849_reg_12434 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_854_fu_6722_p2 = (add_ln703_853_fu_6718_p2 + add_ln703_852_fu_6713_p2);

assign add_ln703_855_fu_6882_p2 = (sub_ln703_759_reg_12525 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_856_fu_6891_p2 = (add_ln703_849_reg_12434_pp0_iter14_reg + sub_ln703_742_fu_6799_p2);

assign add_ln703_857_fu_6728_p2 = (sub_ln703_716_fu_6354_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_858_fu_6733_p2 = (add_ln703_853_fu_6718_p2 + add_ln703_857_fu_6728_p2);

assign add_ln703_859_fu_6901_p2 = (sub_ln703_761_reg_12530 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_860_fu_6905_p2 = (add_ln703_849_reg_12434_pp0_iter14_reg + sub_ln703_745_fu_6807_p2);

assign add_ln703_861_fu_6919_p2 = (sub_ln703_763_reg_12540 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_862_fu_6923_p2 = (sub_ln703_764_fu_6845_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_863_fu_6744_p2 = (add_ln703_816_reg_12241_pp0_iter13_reg + sub_ln703_706_fu_6298_p2);

assign add_ln703_864_fu_6749_p2 = (add_ln703_853_fu_6718_p2 + add_ln703_863_fu_6744_p2);

assign add_ln703_865_fu_6968_p2 = (sub_ln703_770_reg_12570 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_866_fu_6972_p2 = (sub_ln703_724_reg_12450 + data_50_V_read51_reg_8984_pp0_iter14_reg);

assign add_ln703_867_fu_6234_p2 = (data_52_V_read_3_reg_8928_pp0_iter12_reg + data_53_V_read_3_reg_8899_pp0_iter12_reg);

assign add_ln703_868_fu_6755_p2 = (add_ln703_867_reg_12444 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_869_fu_6976_p2 = (add_ln703_868_reg_12585 + add_ln703_866_fu_6972_p2);

assign add_ln703_870_fu_7025_p2 = (sub_ln703_777_fu_6928_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_871_fu_7040_p2 = (sub_ln703_782_fu_6946_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_872_fu_7050_p2 = (sub_ln703_784_fu_6954_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_873_fu_7055_p2 = (sub_ln703_785_fu_6959_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_874_fu_7084_p2 = (sub_ln703_791_fu_6996_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_875_fu_7094_p2 = (sub_ln703_793_fu_7005_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_876_fu_6769_p2 = (add_ln703_826_reg_12419 + sub_ln703_717_fu_6364_p2);

assign add_ln703_877_fu_6774_p2 = (data_53_V_read_3_reg_8899_pp0_iter13_reg + data_54_V_read_3_reg_8873_pp0_iter13_reg);

assign add_ln703_878_fu_7104_p2 = (add_ln703_877_reg_12605 + add_ln703_849_reg_12434_pp0_iter14_reg);

assign add_ln703_879_fu_7108_p2 = (add_ln703_878_fu_7104_p2 + add_ln703_876_reg_12600);

assign add_ln703_880_fu_7113_p2 = (sub_ln703_746_reg_12500 + data_51_V_read52_reg_8956_pp0_iter14_reg);

assign add_ln703_881_fu_7117_p2 = (add_ln703_877_reg_12605 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_882_fu_7121_p2 = (add_ln703_881_fu_7117_p2 + add_ln703_880_fu_7113_p2);

assign add_ln703_883_fu_7127_p2 = (sub_ln703_795_fu_7015_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_884_fu_7132_p2 = (sub_ln703_796_fu_7020_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_885_fu_7142_p2 = (sub_ln703_798_fu_7035_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_886_fu_7147_p2 = (add_ln703_877_reg_12605 + sub_ln703_781_reg_12580);

assign add_ln703_887_fu_7151_p2 = (sub_ln703_768_fu_6858_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_888_fu_7156_p2 = (add_ln703_877_reg_12605 + add_ln703_887_fu_7151_p2);

assign add_ln703_889_fu_7161_p2 = (sub_ln703_799_reg_12595 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_890_fu_7354_p2 = (sub_ln703_801_reg_12660 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_891_fu_7358_p2 = (sub_ln703_802_reg_12665 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_892_fu_7175_p2 = (sub_ln703_803_fu_7070_p2 + data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign add_ln703_893_fu_7180_p2 = (sub_ln703_804_fu_7075_p2 + data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign add_ln703_894_fu_6778_p2 = (data_54_V_read_3_reg_8873_pp0_iter13_reg + data_55_V_read_3_reg_8844_pp0_iter13_reg);

assign add_ln703_895_fu_7185_p2 = (add_ln703_894_reg_12616 + sub_ln703_788_fu_6981_p2);

assign add_ln703_896_fu_7190_p2 = (sub_ln703_773_fu_6886_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_897_fu_7362_p2 = (add_ln703_894_reg_12616_pp0_iter15_reg + add_ln703_896_reg_12725);

assign add_ln703_898_fu_7195_p2 = (sub_ln703_774_fu_6896_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_899_fu_7366_p2 = (add_ln703_894_reg_12616_pp0_iter15_reg + add_ln703_898_reg_12730);

assign add_ln703_900_fu_7378_p2 = (sub_ln703_807_reg_12685 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_901_fu_7390_p2 = (sub_ln703_808_reg_12700 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_902_fu_7394_p2 = (add_ln703_894_reg_12616_pp0_iter15_reg + sub_ln703_797_reg_12645);

assign add_ln703_903_fu_7402_p2 = (sub_ln703_811_fu_7346_p2 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_904_fu_7240_p2 = (sub_ln703_789_fu_6986_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_905_fu_6782_p2 = (data_55_V_read_3_reg_8844_pp0_iter13_reg + data_56_V_read_3_reg_8814_pp0_iter13_reg);

assign add_ln703_906_fu_7245_p2 = (add_ln703_905_reg_12625 + add_ln703_904_fu_7240_p2);

assign add_ln703_907_fu_7477_p2 = (sub_ln703_820_reg_12750 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_908_fu_7250_p2 = (sub_ln703_780_fu_6942_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_909_fu_7255_p2 = (add_ln703_905_reg_12625 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_910_fu_7259_p2 = (add_ln703_909_fu_7255_p2 + add_ln703_908_fu_7250_p2);

assign add_ln703_911_fu_7481_p2 = (sub_ln703_821_reg_12755 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_912_fu_7490_p2 = (sub_ln703_824_reg_12765 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_913_fu_7494_p2 = (sub_ln703_825_reg_12770 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_914_fu_6786_p2 = (sub_ln703_738_fu_6521_p2 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_915_fu_7265_p2 = (add_ln703_849_reg_12434_pp0_iter14_reg + add_ln703_914_reg_12632);

assign add_ln703_916_fu_7269_p2 = (add_ln703_905_reg_12625 + add_ln703_877_reg_12605);

assign add_ln703_917_fu_7273_p2 = (add_ln703_916_fu_7269_p2 + add_ln703_915_fu_7265_p2);

assign add_ln703_918_fu_7513_p2 = (sub_ln703_828_fu_7417_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_919_fu_7279_p2 = (add_ln703_867_reg_12444_pp0_iter14_reg + sub_ln703_757_reg_12515);

assign add_ln703_920_fu_6791_p2 = (data_56_V_read_3_reg_8814_pp0_iter13_reg + data_57_V_read_3_reg_8786_pp0_iter13_reg);

assign add_ln703_921_fu_7283_p2 = (add_ln703_920_reg_12637 + add_ln703_894_reg_12616);

assign add_ln703_922_fu_7287_p2 = (add_ln703_921_fu_7283_p2 + add_ln703_919_fu_7279_p2);

assign add_ln703_923_fu_7293_p2 = (add_ln703_877_reg_12605 + sub_ln703_771_fu_6873_p2);

assign add_ln703_924_fu_7298_p2 = (add_ln703_920_reg_12637 + data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign add_ln703_925_fu_7302_p2 = (add_ln703_924_fu_7298_p2 + add_ln703_923_fu_7293_p2);

assign add_ln703_926_fu_7532_p2 = (sub_ln703_832_fu_7434_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_927_fu_7537_p2 = (sub_ln703_805_reg_12670 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_928_fu_7541_p2 = (add_ln703_920_reg_12637_pp0_iter15_reg + add_ln703_927_fu_7537_p2);

assign add_ln703_929_fu_7546_p2 = (sub_ln703_833_fu_7439_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_930_fu_7561_p2 = (sub_ln703_837_fu_7458_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_931_fu_7308_p2 = (add_ln703_877_reg_12605 + sub_ln703_776_fu_6915_p2);

assign add_ln703_932_fu_7313_p2 = (add_ln703_924_fu_7298_p2 + add_ln703_931_fu_7308_p2);

assign add_ln703_933_fu_7581_p2 = (sub_ln703_841_fu_7485_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_934_fu_7610_p2 = (sub_ln703_844_fu_7508_p2 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_935_fu_7629_p2 = (sub_ln703_846_fu_7523_p2 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_936_fu_7634_p2 = (sub_ln703_847_fu_7528_p2 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_937_fu_7659_p2 = (data_57_V_read_3_reg_8786_pp0_iter15_reg + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_938_fu_7663_p2 = (add_ln703_937_fu_7659_p2 + sub_ln703_835_fu_7449_p2);

assign add_ln703_939_fu_7679_p2 = (add_ln703_937_fu_7659_p2 + sub_ln703_838_fu_7463_p2);

assign add_ln703_940_fu_7690_p2 = (add_ln703_937_fu_7659_p2 + sub_ln703_840_fu_7472_p2);

assign add_ln703_941_fu_7701_p2 = (sub_ln703_852_reg_12790 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_942_fu_7715_p2 = (sub_ln703_823_reg_12760 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_943_fu_7719_p2 = (add_ln703_937_fu_7659_p2 + add_ln703_942_fu_7715_p2);

assign add_ln703_944_fu_7882_p2 = (sub_ln703_858_reg_12840 + data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign add_ln703_945_fu_7740_p2 = (sub_ln703_830_fu_7426_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_946_fu_7334_p2 = (data_58_V_read_3_reg_8756_pp0_iter14_reg + data_59_V_read_3_reg_8724_pp0_iter14_reg);

assign add_ln703_947_fu_7745_p2 = (add_ln703_946_reg_12805 + add_ln703_945_fu_7740_p2);

assign add_ln703_948_fu_7760_p2 = (sub_ln703_864_fu_7644_p2 + data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign add_ln703_949_fu_7765_p2 = (sub_ln703_817_fu_7382_p2 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_950_fu_7770_p2 = (add_ln703_946_reg_12805 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_951_fu_7774_p2 = (add_ln703_950_fu_7770_p2 + add_ln703_949_fu_7765_p2);

assign add_ln703_952_fu_7800_p2 = (add_ln703_946_reg_12805 + sub_ln703_854_fu_7586_p2);

assign add_ln703_953_fu_7956_p2 = (sub_ln703_877_fu_7886_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_954_fu_7338_p2 = (data_59_V_read_3_reg_8724_pp0_iter14_reg + data_60_V_read61_reg_8691_pp0_iter14_reg);

assign add_ln703_955_fu_7815_p2 = (add_ln703_954_reg_12812 + sub_ln703_862_reg_12795);

assign add_ln703_956_fu_7819_p2 = (add_ln703_920_reg_12637_pp0_iter15_reg + sub_ln703_816_reg_12740);

assign add_ln703_957_fu_7823_p2 = (add_ln703_954_reg_12812 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_958_fu_7827_p2 = (add_ln703_957_fu_7823_p2 + add_ln703_956_fu_7819_p2);

assign add_ln703_959_fu_7997_p2 = (sub_ln703_889_fu_7922_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_960_fu_8012_p2 = (sub_ln703_892_reg_12935 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_961_fu_8016_p2 = (sub_ln703_893_reg_12940 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_962_fu_8052_p2 = (sub_ln703_905_fu_7970_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_963_fu_8062_p2 = (sub_ln703_908_fu_7983_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_964_fu_7848_p2 = (data_60_V_read61_reg_8691_pp0_iter15_reg + data_61_V_read62_reg_8663_pp0_iter15_reg);

assign add_ln703_965_fu_8067_p2 = (add_ln703_964_reg_12985 + sub_ln703_886_fu_7910_p2);

assign add_ln703_966_fu_8100_p2 = (sub_ln703_914_fu_8020_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_967_fu_8105_p2 = (sub_ln703_915_fu_8024_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_968_fu_8110_p2 = (add_ln703_964_reg_12985 + sub_ln703_897_fu_7938_p2);

assign add_ln703_969_fu_8115_p2 = (sub_ln703_918_fu_8033_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_970_fu_8125_p2 = (data_61_V_read62_reg_8663_pp0_iter16_reg + data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign add_ln703_971_fu_8129_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_904_reg_12960);

assign add_ln703_972_fu_8148_p2 = (sub_ln703_882_fu_7894_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_973_fu_8153_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_972_fu_8148_p2);

assign add_ln703_974_fu_8159_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_907_fu_7978_p2);

assign add_ln703_975_fu_8170_p2 = (sub_ln703_884_fu_7902_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_976_fu_8175_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_975_fu_8170_p2);

assign add_ln703_977_fu_8186_p2 = (sub_ln703_887_fu_7914_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_978_fu_8191_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_977_fu_8186_p2);

assign add_ln703_979_fu_8197_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_910_fu_7992_p2);

assign add_ln703_980_fu_8203_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_912_fu_8002_p2);

assign add_ln703_981_fu_8214_p2 = (sub_ln703_929_fu_8095_p2 + data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign add_ln703_982_fu_8239_p2 = (sub_ln703_899_fu_7942_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_983_fu_8244_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_982_fu_8239_p2);

assign add_ln703_984_fu_8250_p2 = (sub_ln703_900_fu_7946_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_985_fu_7342_p2 = (data_62_V_read_3_reg_8645_pp0_iter14_reg + data_63_V_read_3_reg_8620_pp0_iter14_reg);

assign add_ln703_986_fu_8255_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_984_fu_8250_p2);

assign add_ln703_987_fu_8260_p2 = (sub_ln703_901_fu_7951_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_994_fu_8325_p2 = (sub_ln703_909_fu_7987_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_fu_530_p2 = (data_0_V_read_int_reg + data_1_V_read_int_reg);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign sub_ln703_100_fu_1329_p2 = (add_ln703_199_fu_1213_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_101_fu_1334_p2 = (sub_ln703_83_fu_1218_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_102_fu_1344_p2 = (add_ln703_200_fu_1226_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_103_fu_1363_p2 = (sub_ln703_87_fu_1238_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_104_fu_1368_p2 = (add_ln703_201_fu_1243_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_105_fu_1373_p2 = (sub_ln703_88_fu_1248_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_106_fu_1378_p2 = (sub_ln703_89_fu_1252_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_107_fu_1383_p2 = (sub_ln703_90_fu_1257_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_108_fu_1388_p2 = (sub_ln703_91_fu_1261_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_109_fu_1407_p2 = (add_ln703_202_fu_1265_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_10_fu_615_p2 = (data_3_V_read_10_reg_10295_pp0_iter2_reg - add_ln703_131_reg_10354_pp0_iter2_reg);

assign sub_ln703_110_fu_1412_p2 = (add_ln703_203_fu_1270_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_111_fu_1417_p2 = (sub_ln703_93_fu_1275_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_112_fu_1422_p2 = (sub_ln703_94_fu_1280_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_113_fu_1427_p2 = (add_ln703_206_fu_1290_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_114_fu_1630_p2 = (add_ln703_207_reg_10682 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_115_fu_1432_p2 = (sub_ln703_97_fu_1304_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_116_fu_1634_p2 = (add_ln703_208_reg_10687 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_117_fu_1638_p2 = (add_ln703_210_reg_10692 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_118_fu_1642_p2 = (sub_ln703_98_reg_10697 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_119_fu_1442_p2 = (sub_ln703_99_fu_1324_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_11_fu_576_p2 = (sub_ln703_5_fu_564_p2 - data_3_V_read_10_reg_10295_pp0_iter1_reg);

assign sub_ln703_120_fu_1447_p2 = (add_ln703_211_fu_1339_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_121_fu_1646_p2 = (add_ln703_216_reg_10702 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_122_fu_1462_p2 = (add_ln703_215_fu_1353_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_123_fu_1467_p2 = (sub_ln703_103_fu_1363_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_124_fu_1650_p2 = (sub_ln703_106_reg_10707 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_125_fu_1482_p2 = (add_ln703_219_fu_1397_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_126_fu_1487_p2 = (add_ln703_221_fu_1402_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_127_fu_1662_p2 = (sub_ln703_109_reg_10722 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_128_fu_1496_p2 = (sub_ln703_111_fu_1417_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_129_fu_1506_p2 = (sub_ln703_113_fu_1427_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_12_fu_627_p2 = (add_ln703_131_reg_10354_pp0_iter2_reg - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_130_fu_1666_p2 = (add_ln703_222_fu_1626_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_131_fu_1680_p2 = (add_ln703_224_reg_10732 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_132_fu_1684_p2 = (sub_ln703_118_fu_1642_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_133_fu_1532_p2 = (add_ln703_225_fu_1452_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_134_fu_1689_p2 = (add_ln703_226_reg_10737 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_135_fu_1698_p2 = (sub_ln703_123_reg_10747 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_136_fu_1702_p2 = (add_ln703_227_reg_10752 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_137_fu_1548_p2 = (add_ln703_228_fu_1477_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_138_fu_1706_p2 = (sub_ln703_124_fu_1650_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_139_fu_1711_p2 = (add_ln703_229_fu_1654_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_13_fu_689_p2 = (sub_ln703_6_reg_10408 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_140_fu_1716_p2 = (add_ln703_230_fu_1658_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_141_fu_1553_p2 = (sub_ln703_126_fu_1487_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_142_fu_1558_p2 = (add_ln703_232_fu_1492_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_143_fu_1725_p2 = (sub_ln703_127_fu_1662_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_144_fu_1730_p2 = (sub_ln703_128_reg_10762 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_145_fu_1734_p2 = (add_ln703_233_reg_10767 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_146_fu_1580_p2 = (sub_ln703_129_fu_1506_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_147_fu_1738_p2 = (sub_ln703_130_fu_1666_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_148_fu_1743_p2 = (add_ln703_234_fu_1671_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_149_fu_1748_p2 = (add_ln703_235_fu_1676_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_14_fu_693_p2 = (add_ln703_132_reg_10414 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_150_fu_1763_p2 = (add_ln703_236_reg_10772 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_151_fu_1767_p2 = (add_ln703_238_reg_10777 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_152_fu_1599_p2 = (add_ln703_240_fu_1526_p2 - data_13_V_read14_reg_10015_pp0_iter4_reg);

assign sub_ln703_153_fu_1775_p2 = (add_ln703_241_fu_1693_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_154_fu_1609_p2 = (add_ln703_244_fu_1542_p2 - data_13_V_read14_reg_10015_pp0_iter4_reg);

assign sub_ln703_155_fu_1780_p2 = (sub_ln703_135_fu_1698_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_156_fu_1785_p2 = (sub_ln703_136_fu_1702_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_157_fu_1790_p2 = (sub_ln703_137_reg_10787 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_158_fu_1794_p2 = (sub_ln703_139_fu_1711_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_159_fu_1799_p2 = (sub_ln703_140_fu_1716_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_15_fu_631_p2 = (add_ln703_133_fu_603_p2 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_160_fu_1804_p2 = (add_ln703_245_fu_1721_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_161_fu_1809_p2 = (sub_ln703_141_reg_10792 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_162_fu_1813_p2 = (sub_ln703_142_reg_10797 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_163_fu_1817_p2 = (add_ln703_247_reg_10802 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_164_fu_1826_p2 = (add_ln703_250_reg_10807 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_165_fu_1830_p2 = (sub_ln703_146_reg_10812 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_166_fu_1834_p2 = (sub_ln703_148_fu_1743_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_167_fu_1839_p2 = (sub_ln703_149_fu_1748_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_168_fu_1844_p2 = (add_ln703_251_fu_1753_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_169_fu_1849_p2 = (add_ln703_253_fu_1758_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_16_fu_640_p2 = (data_4_V_read_10_reg_10273_pp0_iter2_reg - add_ln703_134_reg_10385);

assign sub_ln703_170_fu_1859_p2 = (sub_ln703_150_fu_1763_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_171_fu_1864_p2 = (add_ln703_260_reg_10817 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_172_fu_1868_p2 = (sub_ln703_151_fu_1767_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_173_fu_1873_p2 = (sub_ln703_152_reg_10822 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_174_fu_1877_p2 = (add_ln703_262_reg_10827 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_175_fu_1881_p2 = (add_ln703_263_fu_1771_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_176_fu_1900_p2 = (sub_ln703_154_reg_10832 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_177_fu_1904_p2 = (sub_ln703_156_fu_1785_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_178_fu_1909_p2 = (sub_ln703_157_fu_1790_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_179_fu_1919_p2 = (sub_ln703_160_fu_1804_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_17_fu_653_p2 = (sub_ln703_9_fu_611_p2 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_180_fu_1929_p2 = (sub_ln703_162_fu_1813_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_181_fu_1944_p2 = (add_ln703_264_fu_1821_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_182_fu_1949_p2 = (sub_ln703_164_fu_1826_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_183_fu_1959_p2 = (sub_ln703_168_fu_1844_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_184_fu_1984_p2 = (add_ln703_266_fu_1854_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_185_fu_1989_p2 = (sub_ln703_172_fu_1868_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_186_fu_1994_p2 = (sub_ln703_173_fu_1873_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_187_fu_1999_p2 = (sub_ln703_174_fu_1877_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_188_fu_2004_p2 = (add_ln703_268_fu_1886_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_189_fu_2014_p2 = (add_ln703_271_fu_1895_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_18_fu_658_p2 = (sub_ln703_8_reg_10392 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_190_fu_2024_p2 = (sub_ln703_178_fu_1909_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_191_fu_2029_p2 = (add_ln703_273_fu_1914_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_192_fu_2044_p2 = (add_ln703_274_fu_1924_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_193_fu_2049_p2 = (sub_ln703_180_fu_1929_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_194_fu_2054_p2 = (add_ln703_276_fu_1934_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_195_fu_2059_p2 = (add_ln703_277_fu_1939_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_196_fu_2074_p2 = (sub_ln703_181_fu_1944_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_197_fu_2079_p2 = (add_ln703_278_fu_1954_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_198_fu_2099_p2 = (add_ln703_282_fu_1973_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_199_fu_2246_p2 = (add_ln703_283_reg_10873 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_19_fu_705_p2 = (sub_ln703_10_reg_10420 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_1_fu_540_p2 = (data_0_V_read_10_reg_10329 - data_1_V_read_10_reg_10323);

assign sub_ln703_200_fu_2115_p2 = (sub_ln703_188_fu_2004_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_201_fu_2258_p2 = (add_ln703_285_reg_10888 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_202_fu_2120_p2 = (sub_ln703_189_fu_2014_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_203_fu_2131_p2 = (add_ln703_287_fu_2019_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_204_fu_2142_p2 = (sub_ln703_190_fu_2024_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_205_fu_2262_p2 = (sub_ln703_191_reg_10893 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_206_fu_2266_p2 = (add_ln703_289_reg_10898 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_207_fu_2274_p2 = (add_ln703_290_reg_10903 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_208_fu_2152_p2 = (sub_ln703_192_fu_2044_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_209_fu_2157_p2 = (sub_ln703_195_fu_2059_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_20_fu_662_p2 = (add_ln703_134_reg_10385 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_210_fu_2162_p2 = (add_ln703_293_fu_2069_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_211_fu_2278_p2 = (sub_ln703_196_reg_10913 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_212_fu_2173_p2 = (sub_ln703_197_fu_2079_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_213_fu_2282_p2 = (add_ln703_296_fu_2238_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_214_fu_2287_p2 = (add_ln703_298_fu_2242_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_215_fu_2292_p2 = (add_ln703_300_reg_10930 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_216_fu_2296_p2 = (sub_ln703_198_reg_10935 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_217_fu_2305_p2 = (add_ln703_301_fu_2250_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_218_fu_2310_p2 = (add_ln703_303_reg_10940 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_219_fu_2314_p2 = (add_ln703_304_reg_10945 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_21_fu_709_p2 = (sub_ln703_11_reg_10398_pp0_iter3_reg - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_220_fu_2318_p2 = (add_ln703_305_fu_2254_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_221_fu_2332_p2 = (add_ln703_307_reg_10960 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_222_fu_2340_p2 = (add_ln703_309_reg_10970 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_223_fu_2344_p2 = (sub_ln703_204_reg_10975 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_224_fu_2348_p2 = (sub_ln703_205_fu_2262_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_225_fu_2358_p2 = (add_ln703_312_fu_2270_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_226_fu_2363_p2 = (sub_ln703_207_fu_2274_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_227_fu_2368_p2 = (sub_ln703_209_reg_10990 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_228_fu_2372_p2 = (sub_ln703_210_reg_10995 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_229_fu_2376_p2 = (sub_ln703_211_fu_2278_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_22_fu_713_p2 = (add_ln703_135_reg_10425 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_230_fu_2194_p2 = (add_ln703_314_fu_2167_p2 - data_17_V_read18_reg_9904_pp0_iter5_reg);

assign sub_ln703_231_fu_2381_p2 = (sub_ln703_212_reg_11000 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_232_fu_2385_p2 = (sub_ln703_213_fu_2282_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_233_fu_2390_p2 = (sub_ln703_215_fu_2292_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_234_fu_2395_p2 = (sub_ln703_216_fu_2296_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_235_fu_2400_p2 = (add_ln703_315_fu_2300_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_236_fu_2415_p2 = (sub_ln703_220_fu_2318_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_237_fu_2214_p2 = (add_ln703_317_fu_2182_p2 - data_18_V_read_8_reg_9874_pp0_iter5_reg);

assign sub_ln703_238_fu_2424_p2 = (add_ln703_318_fu_2323_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_239_fu_2429_p2 = (add_ln703_319_fu_2328_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_23_fu_666_p2 = (add_ln703_136_fu_623_p2 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_240_fu_2434_p2 = (sub_ln703_221_fu_2332_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_241_fu_2439_p2 = (add_ln703_320_fu_2336_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_242_fu_2444_p2 = (sub_ln703_222_fu_2340_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_243_fu_2454_p2 = (add_ln703_321_fu_2353_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_244_fu_2468_p2 = (add_ln703_323_reg_11005 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_245_fu_2472_p2 = (sub_ln703_227_fu_2368_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_246_fu_2477_p2 = (sub_ln703_228_fu_2372_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_247_fu_2482_p2 = (sub_ln703_229_fu_2376_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_248_fu_2487_p2 = (sub_ln703_230_reg_11010 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_249_fu_2496_p2 = (sub_ln703_232_fu_2385_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_24_fu_717_p2 = (sub_ln703_13_fu_689_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_250_fu_2501_p2 = (sub_ln703_235_fu_2400_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_251_fu_2506_p2 = (add_ln703_324_fu_2405_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_252_fu_2511_p2 = (add_ln703_328_reg_11015 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_253_fu_2515_p2 = (add_ln703_329_fu_2410_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_254_fu_2525_p2 = (sub_ln703_236_fu_2415_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_255_fu_2530_p2 = (add_ln703_333_reg_11025 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_256_fu_2534_p2 = (add_ln703_335_fu_2420_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_257_fu_2539_p2 = (sub_ln703_238_fu_2424_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_258_fu_2544_p2 = (sub_ln703_239_fu_2429_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_259_fu_2549_p2 = (sub_ln703_240_fu_2434_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_25_fu_722_p2 = (sub_ln703_14_fu_693_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_260_fu_2559_p2 = (sub_ln703_242_fu_2444_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_261_fu_2569_p2 = (add_ln703_336_fu_2449_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_262_fu_2574_p2 = (sub_ln703_243_fu_2454_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_263_fu_2579_p2 = (add_ln703_337_fu_2459_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_264_fu_2584_p2 = (add_ln703_339_fu_2464_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_265_fu_2613_p2 = (sub_ln703_247_fu_2482_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_266_fu_2618_p2 = (sub_ln703_248_fu_2487_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_267_fu_2623_p2 = (add_ln703_340_fu_2491_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_268_fu_2783_p2 = (sub_ln703_249_reg_11056 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_269_fu_2787_p2 = (sub_ln703_251_reg_11066 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_26_fu_727_p2 = (add_ln703_137_fu_697_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_270_fu_2628_p2 = (sub_ln703_252_fu_2511_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_271_fu_2791_p2 = (add_ln703_342_reg_11071 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_272_fu_2647_p2 = (sub_ln703_255_fu_2530_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_273_fu_2799_p2 = (sub_ln703_256_reg_11081 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_274_fu_2652_p2 = (sub_ln703_258_fu_2544_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_275_fu_2662_p2 = (add_ln703_343_fu_2554_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_276_fu_2667_p2 = (add_ln703_345_fu_2564_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_277_fu_2803_p2 = (sub_ln703_261_reg_11091 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_278_fu_2807_p2 = (sub_ln703_262_reg_11096 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_279_fu_2815_p2 = (add_ln703_346_reg_11106 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_27_fu_732_p2 = (sub_ln703_15_reg_10430 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_280_fu_2819_p2 = (add_ln703_350_reg_11111 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_281_fu_2688_p2 = (add_ln703_351_fu_2608_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_282_fu_2827_p2 = (sub_ln703_265_reg_11116 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_283_fu_2693_p2 = (sub_ln703_266_fu_2618_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_284_fu_2698_p2 = (sub_ln703_267_fu_2623_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_285_fu_2836_p2 = (sub_ln703_269_fu_2787_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_286_fu_2845_p2 = (add_ln703_352_reg_11126 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_287_fu_2849_p2 = (sub_ln703_271_fu_2791_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_288_fu_2854_p2 = (add_ln703_353_fu_2795_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_289_fu_2703_p2 = (add_ln703_355_fu_2642_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_28_fu_671_p2 = (data_5_V_read_9_reg_10245_pp0_iter2_reg - add_ln703_139_fu_636_p2);

assign sub_ln703_290_fu_2859_p2 = (sub_ln703_272_reg_11138 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_291_fu_2863_p2 = (sub_ln703_274_reg_11143 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_292_fu_2867_p2 = (add_ln703_356_reg_11148 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_293_fu_2708_p2 = (sub_ln703_276_fu_2667_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_294_fu_2875_p2 = (add_ln703_357_fu_2811_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_295_fu_2880_p2 = (add_ln703_360_reg_11158 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_296_fu_2713_p2 = (add_ln703_361_fu_2683_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_297_fu_2884_p2 = (sub_ln703_279_fu_2815_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_298_fu_2889_p2 = (sub_ln703_280_fu_2819_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_299_fu_2894_p2 = (sub_ln703_281_reg_11163 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_29_fu_749_p2 = (sub_ln703_16_reg_10436 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_2_fu_552_p2 = (sub_ln703_reg_10342 - data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign sub_ln703_300_fu_2898_p2 = (add_ln703_363_fu_2823_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_301_fu_2718_p2 = (sub_ln703_283_fu_2693_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_302_fu_2907_p2 = (add_ln703_364_fu_2831_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_303_fu_2912_p2 = (sub_ln703_285_fu_2836_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_304_fu_2917_p2 = (add_ln703_365_fu_2841_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_305_fu_2922_p2 = (sub_ln703_286_fu_2845_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_306_fu_2931_p2 = (sub_ln703_290_fu_2859_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_307_fu_2941_p2 = (sub_ln703_291_fu_2863_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_308_fu_2946_p2 = (sub_ln703_292_fu_2867_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_309_fu_2951_p2 = (add_ln703_366_fu_2871_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_30_fu_753_p2 = (add_ln703_140_reg_10442 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_310_fu_2978_p2 = (sub_ln703_298_fu_2889_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_311_fu_2988_p2 = (sub_ln703_300_fu_2898_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_312_fu_2993_p2 = (add_ln703_367_fu_2903_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_313_fu_2998_p2 = (sub_ln703_302_fu_2907_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_314_fu_3003_p2 = (add_ln703_371_reg_11193 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_315_fu_3021_p2 = (sub_ln703_303_fu_2912_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_316_fu_3026_p2 = (sub_ln703_304_fu_2917_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_317_fu_3031_p2 = (add_ln703_372_fu_2927_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_318_fu_3036_p2 = (sub_ln703_306_fu_2931_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_319_fu_3041_p2 = (add_ln703_374_fu_2936_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_31_fu_761_p2 = (add_ln703_144_reg_10403_pp0_iter3_reg - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_320_fu_3056_p2 = (sub_ln703_307_fu_2941_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_321_fu_3066_p2 = (sub_ln703_309_fu_2951_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_322_fu_3071_p2 = (add_ln703_377_fu_2956_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_323_fu_3076_p2 = (add_ln703_378_fu_2960_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_324_fu_3091_p2 = (add_ln703_379_fu_2964_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_325_fu_3096_p2 = (add_ln703_380_fu_2969_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_326_fu_3101_p2 = (add_ln703_381_fu_2973_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_327_fu_3106_p2 = (add_ln703_382_fu_2983_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_328_fu_3111_p2 = (sub_ln703_311_fu_2988_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_329_fu_3126_p2 = (sub_ln703_312_fu_2993_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_32_fu_765_p2 = (add_ln703_141_reg_10447 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_330_fu_3372_p2 = (sub_ln703_313_reg_11257 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_331_fu_3140_p2 = (sub_ln703_314_fu_3003_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_332_fu_3376_p2 = (add_ln703_386_reg_11262 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_333_fu_3155_p2 = (sub_ln703_316_fu_3026_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_334_fu_3175_p2 = (sub_ln703_318_fu_3036_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_335_fu_3384_p2 = (add_ln703_390_reg_11272 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_336_fu_3180_p2 = (add_ln703_391_fu_3061_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_337_fu_3190_p2 = (sub_ln703_322_fu_3071_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_338_fu_3195_p2 = (sub_ln703_323_fu_3076_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_339_fu_3200_p2 = (add_ln703_394_fu_3086_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_33_fu_769_p2 = (sub_ln703_18_reg_10459 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_340_fu_3205_p2 = (sub_ln703_324_fu_3091_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_341_fu_3388_p2 = (sub_ln703_326_reg_11277 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_342_fu_3215_p2 = (sub_ln703_327_fu_3106_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_343_fu_3392_p2 = (sub_ln703_328_reg_11282 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_344_fu_3220_p2 = (add_ln703_397_fu_3121_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_345_fu_3234_p2 = (add_ln703_404_fu_3135_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_346_fu_3396_p2 = (add_ln703_410_reg_11287 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_347_fu_3400_p2 = (sub_ln703_332_fu_3376_p2 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_348_fu_3405_p2 = (add_ln703_411_fu_3380_p2 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_349_fu_3410_p2 = (sub_ln703_333_reg_11292 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_34_fu_778_p2 = (sub_ln703_20_reg_10465 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_350_fu_3244_p2 = (add_ln703_413_fu_3160_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_351_fu_3414_p2 = (add_ln703_416_reg_11297 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_352_fu_3427_p2 = (add_ln703_417_reg_11312 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_353_fu_3269_p2 = (sub_ln703_337_fu_3190_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_354_fu_3431_p2 = (sub_ln703_339_reg_11317 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_355_fu_3435_p2 = (sub_ln703_340_reg_11322 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_356_fu_3290_p2 = (add_ln703_418_fu_3210_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_357_fu_3295_p2 = (add_ln703_421_fu_3229_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_358_fu_3300_p2 = (add_ln703_422_fu_3239_p2 - data_26_V_read27_reg_9652_pp0_iter7_reg);

assign sub_ln703_359_fu_3448_p2 = (sub_ln703_349_fu_3410_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_35_fu_787_p2 = (sub_ln703_23_reg_10471 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_360_fu_3453_p2 = (sub_ln703_350_reg_11342 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_361_fu_3457_p2 = (add_ln703_426_reg_11347 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_362_fu_3305_p2 = (add_ln703_428_fu_3264_p2 - data_26_V_read27_reg_9652_pp0_iter7_reg);

assign sub_ln703_363_fu_3461_p2 = (add_ln703_429_fu_3418_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_364_fu_3470_p2 = (add_ln703_430_fu_3423_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_365_fu_3475_p2 = (sub_ln703_352_fu_3427_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_366_fu_3484_p2 = (add_ln703_431_reg_11357 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_367_fu_3488_p2 = (sub_ln703_354_fu_3431_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_368_fu_3493_p2 = (add_ln703_435_reg_11362 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_369_fu_3497_p2 = (sub_ln703_355_fu_3435_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_36_fu_795_p2 = (add_ln703_138_fu_701_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_370_fu_3515_p2 = (add_ln703_436_fu_3439_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_371_fu_3324_p2 = (sub_ln703_357_fu_3295_p2 - data_26_V_read27_reg_9652_pp0_iter7_reg);

assign sub_ln703_372_fu_3532_p2 = (add_ln703_437_fu_3443_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_373_fu_3547_p2 = (sub_ln703_360_fu_3453_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_374_fu_3566_p2 = (add_ln703_440_fu_3466_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_375_fu_3576_p2 = (add_ln703_441_fu_3480_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_376_fu_3591_p2 = (sub_ln703_368_fu_3493_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_377_fu_3596_p2 = (sub_ln703_369_fu_3497_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_378_fu_3601_p2 = (add_ln703_442_fu_3502_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_379_fu_3606_p2 = (add_ln703_444_fu_3506_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_37_fu_800_p2 = (sub_ln703_17_reg_10453 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_380_fu_3611_p2 = (add_ln703_448_fu_3511_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_381_fu_3616_p2 = (sub_ln703_370_fu_3515_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_382_fu_3621_p2 = (add_ln703_450_fu_3520_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_383_fu_3626_p2 = (sub_ln703_371_reg_11397 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_384_fu_3645_p2 = (add_ln703_452_fu_3524_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_385_fu_3650_p2 = (add_ln703_453_fu_3528_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_386_fu_3660_p2 = (add_ln703_455_fu_3537_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_387_fu_3665_p2 = (add_ln703_456_fu_3542_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_388_fu_3670_p2 = (add_ln703_458_fu_3552_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_389_fu_3675_p2 = (add_ln703_461_fu_3561_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_38_fu_814_p2 = (sub_ln703_27_fu_732_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_390_fu_3690_p2 = (add_ln703_462_fu_3571_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_391_fu_3695_p2 = (sub_ln703_375_fu_3576_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_392_fu_3700_p2 = (add_ln703_463_fu_3581_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_393_fu_3705_p2 = (add_ln703_464_fu_3586_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_394_fu_3710_p2 = (sub_ln703_377_fu_3596_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_395_fu_3720_p2 = (sub_ln703_379_fu_3606_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_396_fu_3725_p2 = (sub_ln703_380_fu_3611_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_397_fu_3746_p2 = (sub_ln703_382_fu_3621_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_398_fu_3751_p2 = (sub_ln703_383_fu_3626_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_399_fu_3761_p2 = (add_ln703_468_fu_3639_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_39_fu_819_p2 = (add_ln703_145_fu_736_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_3_fu_560_p2 = (sub_ln703_1_reg_10348 - data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign sub_ln703_400_fu_3973_p2 = (add_ln703_469_reg_11479 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_401_fu_3781_p2 = (sub_ln703_388_fu_3670_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_402_fu_3786_p2 = (sub_ln703_389_fu_3675_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_403_fu_3791_p2 = (add_ln703_474_fu_3680_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_404_fu_3977_p2 = (add_ln703_476_reg_11494 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_405_fu_3816_p2 = (sub_ln703_392_fu_3700_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_406_fu_3981_p2 = (sub_ln703_393_reg_11504 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_407_fu_3985_p2 = (sub_ln703_394_reg_11509 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_408_fu_3845_p2 = (add_ln703_477_fu_3715_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_409_fu_3989_p2 = (sub_ln703_395_reg_11514 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_40_fu_824_p2 = (add_ln703_146_fu_741_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_410_fu_3993_p2 = (add_ln703_478_reg_11519 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_411_fu_3850_p2 = (add_ln703_482_fu_3740_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_412_fu_3855_p2 = (add_ln703_487_fu_3756_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_413_fu_3997_p2 = (sub_ln703_399_reg_11524 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_414_fu_3860_p2 = (add_ln703_488_fu_3766_p2 - data_30_V_read31_reg_9549_pp0_iter8_reg);

assign sub_ln703_415_fu_4001_p2 = (sub_ln703_400_fu_3973_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_416_fu_3865_p2 = (add_ln703_491_fu_3776_p2 - data_30_V_read31_reg_9549_pp0_iter8_reg);

assign sub_ln703_417_fu_4010_p2 = (sub_ln703_402_reg_11534 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_418_fu_4014_p2 = (sub_ln703_404_fu_3977_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_419_fu_3884_p2 = (add_ln703_493_fu_3796_p2 - data_30_V_read31_reg_9549_pp0_iter8_reg);

assign sub_ln703_41_fu_829_p2 = (sub_ln703_28_reg_10476 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_420_fu_4019_p2 = (add_ln703_496_reg_11544 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_421_fu_4023_p2 = (add_ln703_497_reg_11549 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_422_fu_4027_p2 = (sub_ln703_405_reg_11554 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_423_fu_4031_p2 = (add_ln703_506_reg_11559 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_424_fu_4040_p2 = (sub_ln703_408_reg_11564 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_425_fu_4044_p2 = (sub_ln703_409_fu_3989_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_426_fu_4049_p2 = (sub_ln703_410_fu_3993_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_427_fu_4054_p2 = (sub_ln703_411_reg_11569 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_428_fu_4080_p2 = (add_ln703_508_fu_4006_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_429_fu_4102_p2 = (add_ln703_512_reg_11589 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_42_fu_833_p2 = (add_ln703_147_fu_745_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_430_fu_4106_p2 = (sub_ln703_417_fu_4010_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_431_fu_4120_p2 = (sub_ln703_419_reg_11594 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_432_fu_4124_p2 = (sub_ln703_420_fu_4019_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_433_fu_4129_p2 = (sub_ln703_421_fu_4023_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_434_fu_4134_p2 = (sub_ln703_422_fu_4027_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_435_fu_4144_p2 = (add_ln703_513_fu_4035_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_436_fu_4149_p2 = (sub_ln703_424_fu_4040_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_437_fu_4154_p2 = (add_ln703_515_reg_11599 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_438_fu_4163_p2 = (sub_ln703_427_fu_4054_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_439_fu_4168_p2 = (add_ln703_517_reg_11604 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_43_fu_838_p2 = (sub_ln703_29_fu_749_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_440_fu_3938_p2 = (add_ln703_519_fu_3899_p2 - data_31_V_read32_reg_9521_pp0_iter8_reg);

assign sub_ln703_441_fu_4172_p2 = (add_ln703_520_fu_4058_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_442_fu_4177_p2 = (add_ln703_521_fu_4062_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_443_fu_4182_p2 = (add_ln703_522_fu_4067_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_444_fu_4187_p2 = (add_ln703_538_fu_4075_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_445_fu_4192_p2 = (sub_ln703_428_fu_4080_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_446_fu_4197_p2 = (add_ln703_541_fu_4089_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_447_fu_4202_p2 = (add_ln703_545_reg_11614 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_448_fu_4206_p2 = (add_ln703_546_fu_4094_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_449_fu_4211_p2 = (add_ln703_548_fu_4098_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_44_fu_848_p2 = (add_ln703_148_fu_757_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_450_fu_4221_p2 = (sub_ln703_430_fu_4106_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_451_fu_4226_p2 = (add_ln703_550_fu_4111_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_452_fu_4231_p2 = (add_ln703_551_fu_4115_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_453_fu_4236_p2 = (sub_ln703_431_fu_4120_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_454_fu_4246_p2 = (add_ln703_552_fu_4139_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_455_fu_4251_p2 = (add_ln703_556_reg_11619 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_456_fu_4255_p2 = (sub_ln703_436_fu_4149_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_457_fu_4265_p2 = (sub_ln703_437_fu_4154_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_458_fu_4270_p2 = (add_ln703_557_fu_4158_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_459_fu_4284_p2 = (sub_ln703_441_fu_4172_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_45_fu_853_p2 = (sub_ln703_31_fu_761_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_460_fu_4289_p2 = (sub_ln703_443_fu_4182_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_461_fu_4303_p2 = (sub_ln703_445_fu_4192_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_462_fu_4313_p2 = (sub_ln703_447_fu_4202_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_463_fu_4558_p2 = (sub_ln703_448_reg_11673 - data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign sub_ln703_464_fu_4318_p2 = (add_ln703_558_fu_4216_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_465_fu_4328_p2 = (sub_ln703_451_fu_4226_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_466_fu_4562_p2 = (sub_ln703_452_reg_11678 - data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign sub_ln703_467_fu_4333_p2 = (add_ln703_559_fu_4241_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_468_fu_4353_p2 = (sub_ln703_454_fu_4246_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_469_fu_4368_p2 = (sub_ln703_456_fu_4255_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_46_fu_858_p2 = (sub_ln703_32_fu_765_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_470_fu_4373_p2 = (add_ln703_561_fu_4260_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_471_fu_4378_p2 = (sub_ln703_457_fu_4265_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_472_fu_4570_p2 = (sub_ln703_458_reg_11688 - data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign sub_ln703_473_fu_4388_p2 = (add_ln703_562_fu_4275_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_474_fu_4393_p2 = (add_ln703_563_fu_4280_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_475_fu_4418_p2 = (add_ln703_571_fu_4298_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_476_fu_4574_p2 = (sub_ln703_461_reg_11693 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_477_fu_4578_p2 = (add_ln703_572_reg_11698 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_478_fu_4582_p2 = (sub_ln703_462_reg_11703 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_479_fu_4586_p2 = (add_ln703_573_reg_11708 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_47_fu_863_p2 = (sub_ln703_33_fu_769_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_480_fu_4590_p2 = (add_ln703_574_fu_4566_p2 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_481_fu_4595_p2 = (sub_ln703_467_reg_11713 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_482_fu_4447_p2 = (add_ln703_576_fu_4338_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_483_fu_4452_p2 = (add_ln703_580_fu_4348_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_484_fu_4599_p2 = (sub_ln703_468_reg_11718 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_485_fu_4603_p2 = (add_ln703_581_reg_11723 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_486_fu_4607_p2 = (add_ln703_583_reg_11728 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_487_fu_4611_p2 = (sub_ln703_470_reg_11738 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_488_fu_4457_p2 = (sub_ln703_471_fu_4378_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_489_fu_4615_p2 = (sub_ln703_472_fu_4570_p2 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_48_fu_877_p2 = (add_ln703_149_fu_773_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_490_fu_4462_p2 = (add_ln703_585_fu_4383_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_491_fu_4467_p2 = (sub_ln703_473_fu_4388_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_492_fu_4472_p2 = (sub_ln703_474_fu_4393_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_493_fu_4624_p2 = (add_ln703_586_reg_11743 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_494_fu_4632_p2 = (add_ln703_590_reg_11748 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_495_fu_4636_p2 = (sub_ln703_475_reg_11753 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_496_fu_4650_p2 = (add_ln703_591_reg_11758 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_497_fu_4654_p2 = (sub_ln703_479_fu_4586_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_498_fu_4659_p2 = (add_ln703_592_reg_11763 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_499_fu_4663_p2 = (sub_ln703_480_fu_4590_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_49_fu_882_p2 = (sub_ln703_34_fu_778_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_4_fu_548_p2 = (add_ln703_reg_10335 - data_2_V_read_10_reg_10312);

assign sub_ln703_500_fu_4668_p2 = (add_ln703_598_reg_11768 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_501_fu_4672_p2 = (sub_ln703_481_fu_4595_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_502_fu_4682_p2 = (sub_ln703_485_fu_4603_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_503_fu_4516_p2 = (sub_ln703_492_fu_4472_p2 - data_35_V_read_3_reg_9410_pp0_iter9_reg);

assign sub_ln703_504_fu_4700_p2 = (add_ln703_601_fu_4620_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_505_fu_4521_p2 = (add_ln703_608_fu_4495_p2 - data_36_V_read_3_reg_9383_pp0_iter9_reg);

assign sub_ln703_506_fu_4705_p2 = (sub_ln703_493_fu_4624_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_507_fu_4710_p2 = (add_ln703_611_fu_4628_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_508_fu_4715_p2 = (sub_ln703_494_fu_4632_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_509_fu_4725_p2 = (add_ln703_612_fu_4640_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_50_fu_887_p2 = (add_ln703_150_fu_782_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_510_fu_4730_p2 = (add_ln703_613_fu_4645_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_511_fu_4735_p2 = (add_ln703_616_reg_11808 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_512_fu_4744_p2 = (sub_ln703_497_fu_4654_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_513_fu_4749_p2 = (sub_ln703_498_fu_4659_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_514_fu_4764_p2 = (sub_ln703_500_fu_4668_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_515_fu_4778_p2 = (add_ln703_617_fu_4677_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_516_fu_4783_p2 = (sub_ln703_502_fu_4682_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_517_fu_4788_p2 = (add_ln703_618_fu_4687_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_518_fu_4798_p2 = (add_ln703_619_fu_4692_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_519_fu_4808_p2 = (add_ln703_620_fu_4696_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_51_fu_897_p2 = (add_ln703_151_fu_791_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_520_fu_4813_p2 = (sub_ln703_503_reg_11813 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_521_fu_4830_p2 = (sub_ln703_506_fu_4705_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_522_fu_4840_p2 = (sub_ln703_508_fu_4715_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_523_fu_4845_p2 = (add_ln703_622_fu_4720_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_524_fu_4850_p2 = (sub_ln703_511_fu_4735_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_525_fu_4855_p2 = (add_ln703_623_fu_4739_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_526_fu_4860_p2 = (sub_ln703_512_fu_4744_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_527_fu_4865_p2 = (add_ln703_626_fu_4759_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_528_fu_4875_p2 = (sub_ln703_514_fu_4764_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_529_fu_4880_p2 = (add_ln703_627_fu_4769_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_52_fu_907_p2 = (sub_ln703_37_fu_800_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_530_fu_4885_p2 = (add_ln703_629_fu_4774_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_531_fu_4890_p2 = (add_ln703_634_reg_11828 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_532_fu_4894_p2 = (sub_ln703_515_fu_4778_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_533_fu_4904_p2 = (sub_ln703_517_fu_4788_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_534_fu_4909_p2 = (add_ln703_636_fu_4793_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_535_fu_4919_p2 = (add_ln703_638_fu_4803_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_536_fu_4924_p2 = (sub_ln703_520_fu_4813_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_537_fu_4929_p2 = (add_ln703_642_fu_4817_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_538_fu_4934_p2 = (add_ln703_643_fu_4821_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_539_fu_4939_p2 = (add_ln703_644_fu_4826_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_53_fu_912_p2 = (add_ln703_152_fu_804_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_540_fu_4944_p2 = (add_ln703_645_fu_4835_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_541_fu_4949_p2 = (sub_ln703_522_fu_4840_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_542_fu_4954_p2 = (sub_ln703_523_fu_4845_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_543_fu_4979_p2 = (sub_ln703_524_fu_4850_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_544_fu_4984_p2 = (sub_ln703_525_fu_4855_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_545_fu_5138_p2 = (sub_ln703_526_reg_11864 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_546_fu_5142_p2 = (sub_ln703_527_reg_11869 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_547_fu_5146_p2 = (add_ln703_647_reg_11874 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_548_fu_5154_p2 = (sub_ln703_532_reg_11884 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_549_fu_5158_p2 = (add_ln703_648_reg_11889 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_54_fu_1086_p2 = (add_ln703_153_reg_10503 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_550_fu_5162_p2 = (sub_ln703_533_reg_11894 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_551_fu_5004_p2 = (add_ln703_649_fu_4914_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_552_fu_5170_p2 = (sub_ln703_539_reg_11909 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_553_fu_5174_p2 = (sub_ln703_540_reg_11914 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_554_fu_5178_p2 = (sub_ln703_542_reg_11924 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_555_fu_5182_p2 = (add_ln703_651_reg_11929 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_556_fu_5024_p2 = (add_ln703_656_fu_4973_p2 - data_39_V_read_3_reg_9301_pp0_iter10_reg);

assign sub_ln703_557_fu_5029_p2 = (sub_ln703_543_fu_4979_p2 - data_39_V_read_3_reg_9301_pp0_iter10_reg);

assign sub_ln703_558_fu_5034_p2 = (add_ln703_658_fu_4989_p2 - data_39_V_read_3_reg_9301_pp0_iter10_reg);

assign sub_ln703_559_fu_5190_p2 = (sub_ln703_546_fu_5142_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_55_fu_1090_p2 = (sub_ln703_38_reg_10508 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_560_fu_5195_p2 = (sub_ln703_547_fu_5146_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_561_fu_5200_p2 = (add_ln703_659_fu_5150_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_562_fu_5205_p2 = (add_ln703_660_reg_11939 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_563_fu_5209_p2 = (sub_ln703_548_fu_5154_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_564_fu_5214_p2 = (sub_ln703_550_fu_5162_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_565_fu_5219_p2 = (add_ln703_661_reg_11944 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_566_fu_5223_p2 = (sub_ln703_551_reg_11949 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_567_fu_5227_p2 = (add_ln703_662_fu_5166_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_568_fu_5232_p2 = (add_ln703_666_reg_11954 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_569_fu_5236_p2 = (add_ln703_668_reg_11959 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_56_fu_1094_p2 = (sub_ln703_39_reg_10513 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_570_fu_5263_p2 = (sub_ln703_557_reg_11969 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_571_fu_5267_p2 = (add_ln703_669_fu_5186_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_572_fu_5276_p2 = (sub_ln703_560_fu_5195_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_573_fu_5101_p2 = (add_ln703_671_fu_5039_p2 - data_40_V_read41_reg_9272_pp0_iter10_reg);

assign sub_ln703_574_fu_5290_p2 = (sub_ln703_562_fu_5205_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_575_fu_5295_p2 = (add_ln703_676_reg_11979 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_576_fu_5299_p2 = (sub_ln703_564_fu_5214_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_577_fu_5304_p2 = (add_ln703_682_reg_11984 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_578_fu_5308_p2 = (sub_ln703_565_fu_5219_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_579_fu_5318_p2 = (sub_ln703_567_fu_5227_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_57_fu_1102_p2 = (sub_ln703_40_reg_10519 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_580_fu_5323_p2 = (sub_ln703_568_fu_5232_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_581_fu_5328_p2 = (add_ln703_685_reg_11989 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_582_fu_5106_p2 = (add_ln703_687_fu_5082_p2 - data_40_V_read41_reg_9272_pp0_iter10_reg);

assign sub_ln703_583_fu_5111_p2 = (add_ln703_689_fu_5087_p2 - data_40_V_read41_reg_9272_pp0_iter10_reg);

assign sub_ln703_584_fu_5341_p2 = (sub_ln703_569_fu_5236_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_585_fu_5346_p2 = (add_ln703_690_fu_5240_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_586_fu_5351_p2 = (add_ln703_692_fu_5245_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_587_fu_5356_p2 = (add_ln703_693_fu_5249_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_588_fu_5370_p2 = (add_ln703_694_fu_5254_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_589_fu_5375_p2 = (add_ln703_695_fu_5259_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_58_fu_922_p2 = (sub_ln703_41_fu_829_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_590_fu_5380_p2 = (sub_ln703_570_fu_5263_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_591_fu_5385_p2 = (sub_ln703_571_fu_5267_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_592_fu_5400_p2 = (add_ln703_696_fu_5272_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_593_fu_5410_p2 = (sub_ln703_572_fu_5276_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_594_fu_5415_p2 = (add_ln703_699_fu_5281_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_595_fu_5420_p2 = (add_ln703_700_fu_5285_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_596_fu_5444_p2 = (sub_ln703_577_fu_5304_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_597_fu_5449_p2 = (add_ln703_701_fu_5313_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_598_fu_5454_p2 = (sub_ln703_579_fu_5318_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_599_fu_5459_p2 = (sub_ln703_580_fu_5323_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_59_fu_1106_p2 = (sub_ln703_43_reg_10524 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_5_fu_564_p2 = (data_2_V_read_10_reg_10312_pp0_iter1_reg - add_ln703_reg_10335_pp0_iter1_reg);

assign sub_ln703_600_fu_5464_p2 = (sub_ln703_581_fu_5328_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_601_fu_5473_p2 = (sub_ln703_583_reg_12017 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_602_fu_5688_p2 = (add_ln703_704_reg_12056 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_603_fu_5491_p2 = (sub_ln703_587_fu_5356_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_604_fu_5496_p2 = (add_ln703_709_fu_5365_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_605_fu_5501_p2 = (sub_ln703_588_fu_5370_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_606_fu_5696_p2 = (sub_ln703_589_reg_12066 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_607_fu_5506_p2 = (sub_ln703_590_fu_5380_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_608_fu_5511_p2 = (sub_ln703_591_fu_5385_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_609_fu_5516_p2 = (add_ln703_712_fu_5395_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_60_fu_927_p2 = (add_ln703_154_fu_843_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_610_fu_5521_p2 = (add_ln703_714_fu_5405_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_611_fu_5704_p2 = (sub_ln703_594_reg_12076 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_612_fu_5526_p2 = (add_ln703_715_fu_5425_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_613_fu_5531_p2 = (add_ln703_716_fu_5429_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_614_fu_5536_p2 = (add_ln703_718_fu_5434_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_615_fu_5708_p2 = (add_ln703_719_reg_12086 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_616_fu_5712_p2 = (sub_ln703_598_reg_12091 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_617_fu_5561_p2 = (sub_ln703_600_fu_5464_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_618_fu_5566_p2 = (add_ln703_720_fu_5469_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_619_fu_5716_p2 = (sub_ln703_602_fu_5688_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_61_fu_932_p2 = (sub_ln703_44_fu_848_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_620_fu_5721_p2 = (add_ln703_721_fu_5692_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_621_fu_5726_p2 = (add_ln703_728_reg_12096 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_622_fu_5730_p2 = (sub_ln703_603_reg_12101 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_623_fu_5734_p2 = (sub_ln703_604_reg_12106 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_624_fu_5596_p2 = (sub_ln703_607_fu_5506_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_625_fu_5742_p2 = (sub_ln703_609_reg_12121 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_626_fu_5746_p2 = (sub_ln703_610_reg_12126 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_627_fu_5750_p2 = (add_ln703_729_fu_5700_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_628_fu_5755_p2 = (sub_ln703_613_reg_12136 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_629_fu_5763_p2 = (sub_ln703_615_fu_5708_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_62_fu_942_p2 = (add_ln703_156_fu_872_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_630_fu_5627_p2 = (add_ln703_730_fu_5541_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_631_fu_5632_p2 = (add_ln703_732_fu_5546_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_632_fu_5768_p2 = (add_ln703_733_reg_12146 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_633_fu_5772_p2 = (add_ln703_734_reg_12151 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_634_fu_5637_p2 = (sub_ln703_617_fu_5561_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_635_fu_5780_p2 = (add_ln703_735_reg_12161 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_636_fu_5784_p2 = (sub_ln703_619_fu_5716_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_637_fu_5642_p2 = (add_ln703_739_fu_5585_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_638_fu_5647_p2 = (add_ln703_741_fu_5591_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_639_fu_5789_p2 = (sub_ln703_620_fu_5721_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_63_fu_947_p2 = (sub_ln703_48_fu_877_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_640_fu_5794_p2 = (sub_ln703_622_fu_5730_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_641_fu_5799_p2 = (sub_ln703_623_fu_5734_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_642_fu_5804_p2 = (add_ln703_742_fu_5738_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_643_fu_5822_p2 = (sub_ln703_625_fu_5742_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_644_fu_5656_p2 = (add_ln703_744_fu_5601_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_645_fu_5827_p2 = (sub_ln703_626_fu_5746_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_646_fu_5832_p2 = (sub_ln703_627_fu_5750_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_647_fu_5846_p2 = (sub_ln703_628_fu_5755_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_648_fu_5661_p2 = (add_ln703_747_fu_5611_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_649_fu_5851_p2 = (add_ln703_748_fu_5759_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_64_fu_957_p2 = (sub_ln703_49_fu_882_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_650_fu_5666_p2 = (add_ln703_753_fu_5621_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_651_fu_5856_p2 = (sub_ln703_629_fu_5763_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_652_fu_5865_p2 = (sub_ln703_632_fu_5768_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_653_fu_5870_p2 = (sub_ln703_633_fu_5772_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_654_fu_5875_p2 = (sub_ln703_634_reg_12181 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_655_fu_5879_p2 = (add_ln703_754_fu_5776_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_656_fu_5884_p2 = (sub_ln703_635_fu_5780_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_657_fu_5889_p2 = (sub_ln703_638_reg_12191 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_658_fu_5898_p2 = (sub_ln703_640_fu_5794_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_659_fu_5903_p2 = (sub_ln703_642_fu_5804_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_65_fu_1110_p2 = (add_ln703_157_reg_10529 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_660_fu_5908_p2 = (add_ln703_756_fu_5809_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_661_fu_5913_p2 = (add_ln703_757_fu_5814_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_662_fu_5918_p2 = (add_ln703_759_fu_5818_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_663_fu_5923_p2 = (sub_ln703_643_fu_5822_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_664_fu_5928_p2 = (sub_ln703_644_reg_12204 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_665_fu_5932_p2 = (sub_ln703_646_fu_5832_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_666_fu_5937_p2 = (add_ln703_761_fu_5837_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_667_fu_5956_p2 = (add_ln703_763_fu_5842_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_668_fu_5971_p2 = (sub_ln703_650_reg_12214 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_669_fu_5975_p2 = (sub_ln703_651_fu_5856_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_66_fu_987_p2 = (add_ln703_160_fu_902_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_670_fu_5980_p2 = (add_ln703_764_fu_5861_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_671_fu_5989_p2 = (sub_ln703_652_fu_5865_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_672_fu_6004_p2 = (sub_ln703_653_fu_5870_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_673_fu_6009_p2 = (sub_ln703_654_fu_5875_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_674_fu_6014_p2 = (sub_ln703_655_fu_5879_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_675_fu_6019_p2 = (sub_ln703_656_fu_5884_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_676_fu_6033_p2 = (sub_ln703_657_fu_5889_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_677_fu_6047_p2 = (add_ln703_766_fu_5893_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_678_fu_6052_p2 = (sub_ln703_658_fu_5898_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_679_fu_6057_p2 = (sub_ln703_659_fu_5903_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_67_fu_1119_p2 = (add_ln703_162_reg_10539 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_680_fu_6062_p2 = (sub_ln703_660_fu_5908_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_681_fu_6238_p2 = (sub_ln703_662_reg_12248 - data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign sub_ln703_682_fu_6067_p2 = (sub_ln703_664_fu_5928_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_683_fu_6242_p2 = (sub_ln703_665_reg_12253 - data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign sub_ln703_684_fu_6072_p2 = (sub_ln703_666_fu_5937_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_685_fu_6246_p2 = (add_ln703_770_reg_12258 - data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign sub_ln703_686_fu_6077_p2 = (add_ln703_771_fu_5961_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_687_fu_6086_p2 = (add_ln703_772_fu_5966_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_688_fu_6091_p2 = (sub_ln703_668_fu_5971_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_689_fu_6096_p2 = (sub_ln703_670_fu_5980_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_68_fu_1133_p2 = (add_ln703_163_fu_1098_p2 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_690_fu_6101_p2 = (add_ln703_774_fu_5985_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_691_fu_6106_p2 = (sub_ln703_671_fu_5989_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_692_fu_6111_p2 = (add_ln703_777_fu_5999_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_693_fu_6116_p2 = (sub_ln703_672_fu_6004_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_694_fu_6126_p2 = (sub_ln703_674_fu_6014_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_695_fu_6254_p2 = (add_ln703_779_reg_12273 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_696_fu_6136_p2 = (add_ln703_781_fu_6029_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_697_fu_6141_p2 = (add_ln703_786_fu_6042_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_698_fu_6267_p2 = (sub_ln703_682_reg_12298 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_699_fu_6271_p2 = (sub_ln703_683_fu_6242_p2 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_69_fu_1138_p2 = (sub_ln703_57_fu_1102_p2 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_6_fu_595_p2 = (sub_ln703_2_reg_10367 - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_700_fu_6172_p2 = (add_ln703_788_fu_6082_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_701_fu_6281_p2 = (sub_ln703_687_reg_12313 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_702_fu_6285_p2 = (sub_ln703_688_reg_12318 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_703_fu_6289_p2 = (add_ln703_789_fu_6250_p2 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_704_fu_6177_p2 = (sub_ln703_689_fu_6096_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_705_fu_6294_p2 = (sub_ln703_691_reg_12328 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_706_fu_6298_p2 = (sub_ln703_693_reg_12338 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_707_fu_6182_p2 = (add_ln703_790_fu_6121_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_708_fu_6302_p2 = (add_ln703_791_reg_12348 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_709_fu_6306_p2 = (sub_ln703_695_fu_6254_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_70_fu_992_p2 = (sub_ln703_60_fu_927_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_710_fu_6311_p2 = (sub_ln703_696_reg_12353 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_711_fu_6328_p2 = (add_ln703_792_reg_12363 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_712_fu_6332_p2 = (add_ln703_793_fu_6258_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_713_fu_6337_p2 = (add_ln703_796_reg_12368 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_714_fu_6345_p2 = (add_ln703_797_fu_6262_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_715_fu_6350_p2 = (add_ln703_798_reg_12373 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_716_fu_6354_p2 = (sub_ln703_698_fu_6267_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_717_fu_6364_p2 = (add_ln703_799_fu_6276_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_718_fu_6382_p2 = (sub_ln703_700_reg_12378 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_719_fu_6386_p2 = (sub_ln703_701_fu_6281_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_71_fu_1002_p2 = (add_ln703_164_fu_937_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_720_fu_6391_p2 = (sub_ln703_702_fu_6285_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_721_fu_6413_p2 = (sub_ln703_707_reg_12388 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_722_fu_6422_p2 = (sub_ln703_709_fu_6306_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_723_fu_6427_p2 = (add_ln703_800_fu_6315_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_724_fu_6432_p2 = (add_ln703_804_fu_6323_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_725_fu_6437_p2 = (sub_ln703_713_fu_6337_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_726_fu_6442_p2 = (add_ln703_805_fu_6341_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_727_fu_6452_p2 = (sub_ln703_715_fu_6350_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_728_fu_6457_p2 = (add_ln703_806_fu_6359_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_729_fu_6462_p2 = (add_ln703_808_fu_6373_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_72_fu_1147_p2 = (sub_ln703_63_reg_10555 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_730_fu_6467_p2 = (add_ln703_809_fu_6378_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_731_fu_6472_p2 = (sub_ln703_718_fu_6382_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_732_fu_6477_p2 = (sub_ln703_719_fu_6386_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_733_fu_6487_p2 = (add_ln703_810_fu_6396_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_734_fu_6492_p2 = (add_ln703_811_fu_6401_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_735_fu_6497_p2 = (add_ln703_812_fu_6405_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_736_fu_6502_p2 = (add_ln703_813_fu_6409_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_737_fu_6507_p2 = (sub_ln703_721_fu_6413_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_738_fu_6521_p2 = (add_ln703_814_fu_6417_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_739_fu_6541_p2 = (sub_ln703_725_fu_6437_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_73_fu_1026_p2 = (add_ln703_165_fu_952_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_740_fu_6560_p2 = (sub_ln703_726_fu_6442_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_741_fu_6795_p2 = (add_ln703_818_reg_12409_pp0_iter14_reg - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_742_fu_6799_p2 = (add_ln703_819_reg_12455 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_743_fu_6803_p2 = (sub_ln703_727_reg_12460 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_744_fu_6565_p2 = (add_ln703_821_reg_12414 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_745_fu_6807_p2 = (sub_ln703_728_reg_12465 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_746_fu_6579_p2 = (sub_ln703_729_fu_6462_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_747_fu_6584_p2 = (sub_ln703_730_fu_6467_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_748_fu_6589_p2 = (sub_ln703_731_fu_6472_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_749_fu_6599_p2 = (add_ln703_822_fu_6482_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_74_fu_1151_p2 = (sub_ln703_64_reg_10560 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_750_fu_6811_p2 = (sub_ln703_733_reg_12470 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_751_fu_6604_p2 = (sub_ln703_734_fu_6492_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_752_fu_6609_p2 = (sub_ln703_735_fu_6497_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_753_fu_6614_p2 = (sub_ln703_737_fu_6507_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_754_fu_6619_p2 = (add_ln703_824_fu_6516_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_755_fu_6819_p2 = (add_ln703_825_reg_12480 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_756_fu_6823_p2 = (add_ln703_827_reg_12485 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_757_fu_6629_p2 = (add_ln703_828_fu_6536_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_758_fu_6827_p2 = (add_ln703_831_reg_12490 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_759_fu_6639_p2 = (sub_ln703_740_fu_6560_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_75_fu_1031_p2 = (add_ln703_168_fu_967_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_760_fu_6831_p2 = (sub_ln703_741_fu_6795_p2 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_761_fu_6644_p2 = (sub_ln703_744_fu_6565_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_762_fu_6841_p2 = (add_ln703_833_reg_12495 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_763_fu_6654_p2 = (sub_ln703_748_fu_6589_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_764_fu_6845_p2 = (add_ln703_834_reg_12505 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_765_fu_6849_p2 = (sub_ln703_749_reg_12510 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_766_fu_6853_p2 = (sub_ln703_750_fu_6811_p2 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_767_fu_6659_p2 = (sub_ln703_751_fu_6604_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_768_fu_6858_p2 = (add_ln703_835_fu_6815_p2 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_769_fu_6684_p2 = (sub_ln703_753_fu_6614_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_76_fu_1155_p2 = (add_ln703_170_reg_10566 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_770_fu_6708_p2 = (add_ln703_837_fu_6624_p2 - data_52_V_read_3_reg_8928_pp0_iter13_reg);

assign sub_ln703_771_fu_6873_p2 = (add_ln703_838_reg_12520 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_772_fu_6877_p2 = (sub_ln703_758_fu_6827_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_773_fu_6886_p2 = (sub_ln703_760_fu_6831_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_774_fu_6896_p2 = (add_ln703_839_fu_6836_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_775_fu_6910_p2 = (sub_ln703_762_fu_6841_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_776_fu_6915_p2 = (add_ln703_840_reg_12535 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_777_fu_6928_p2 = (sub_ln703_765_fu_6849_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_778_fu_6933_p2 = (sub_ln703_766_fu_6853_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_779_fu_6938_p2 = (sub_ln703_767_reg_12545 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_77_fu_1159_p2 = (sub_ln703_65_fu_1110_p2 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_780_fu_6942_p2 = (add_ln703_841_reg_12550 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_781_fu_6739_p2 = (add_ln703_844_fu_6678_p2 - data_52_V_read_3_reg_8928_pp0_iter13_reg);

assign sub_ln703_782_fu_6946_p2 = (sub_ln703_769_reg_12555 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_783_fu_6950_p2 = (add_ln703_845_reg_12560 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_784_fu_6954_p2 = (add_ln703_846_fu_6863_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_785_fu_6959_p2 = (add_ln703_847_fu_6868_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_786_fu_6964_p2 = (add_ln703_851_reg_12565 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_787_fu_6759_p2 = (add_ln703_854_fu_6722_p2 - data_53_V_read_3_reg_8899_pp0_iter13_reg);

assign sub_ln703_788_fu_6981_p2 = (sub_ln703_772_fu_6877_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_789_fu_6986_p2 = (add_ln703_855_fu_6882_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_78_fu_1164_p2 = (add_ln703_171_reg_10571 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_790_fu_6991_p2 = (add_ln703_856_fu_6891_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_791_fu_6996_p2 = (add_ln703_858_reg_12575 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_792_fu_7000_p2 = (add_ln703_859_fu_6901_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_793_fu_7005_p2 = (add_ln703_860_fu_6905_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_794_fu_7010_p2 = (sub_ln703_775_fu_6910_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_795_fu_7015_p2 = (add_ln703_861_fu_6919_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_796_fu_7020_p2 = (add_ln703_862_fu_6923_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_797_fu_7030_p2 = (sub_ln703_778_fu_6933_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_798_fu_7035_p2 = (sub_ln703_779_fu_6938_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_799_fu_6764_p2 = (add_ln703_864_fu_6749_p2 - data_53_V_read_3_reg_8899_pp0_iter13_reg);

assign sub_ln703_79_fu_1168_p2 = (add_ln703_173_reg_10576 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_7_fu_607_p2 = (add_ln703_130_reg_10373 - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_800_fu_7045_p2 = (sub_ln703_783_fu_6950_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_801_fu_7060_p2 = (sub_ln703_786_fu_6964_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_802_fu_7065_p2 = (add_ln703_865_fu_6968_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_803_fu_7070_p2 = (add_ln703_869_fu_6976_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_804_fu_7075_p2 = (sub_ln703_787_reg_12590 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_805_fu_7079_p2 = (sub_ln703_790_fu_6991_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_806_fu_7089_p2 = (sub_ln703_792_fu_7000_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_807_fu_7099_p2 = (sub_ln703_794_fu_7010_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_808_fu_7137_p2 = (add_ln703_870_fu_7025_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_809_fu_7165_p2 = (add_ln703_871_fu_7040_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_80_fu_1184_p2 = (add_ln703_174_fu_1114_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_810_fu_7170_p2 = (sub_ln703_800_fu_7045_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_811_fu_7346_p2 = (add_ln703_872_reg_12650 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_812_fu_7350_p2 = (add_ln703_873_reg_12655 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_813_fu_7370_p2 = (add_ln703_874_reg_12675 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_814_fu_7200_p2 = (sub_ln703_806_fu_7089_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_815_fu_7374_p2 = (add_ln703_875_reg_12680 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_816_fu_7205_p2 = (add_ln703_879_fu_7108_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_817_fu_7382_p2 = (add_ln703_882_reg_12690 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_818_fu_7210_p2 = (add_ln703_883_fu_7127_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_819_fu_7386_p2 = (add_ln703_884_reg_12695 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_81_fu_1194_p2 = (add_ln703_175_fu_1123_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_820_fu_7215_p2 = (add_ln703_885_fu_7142_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_821_fu_7220_p2 = (add_ln703_886_fu_7147_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_822_fu_7398_p2 = (add_ln703_888_reg_12705 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_823_fu_7225_p2 = (add_ln703_889_fu_7161_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_824_fu_7230_p2 = (sub_ln703_809_fu_7165_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_825_fu_7235_p2 = (sub_ln703_810_fu_7170_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_826_fu_7407_p2 = (sub_ln703_812_fu_7350_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_827_fu_7412_p2 = (add_ln703_890_fu_7354_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_828_fu_7417_p2 = (add_ln703_891_fu_7358_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_829_fu_7422_p2 = (add_ln703_892_reg_12710 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_82_fu_1199_p2 = (add_ln703_176_fu_1128_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_830_fu_7426_p2 = (add_ln703_893_reg_12715 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_831_fu_7430_p2 = (add_ln703_895_reg_12720 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_832_fu_7434_p2 = (add_ln703_897_fu_7362_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_833_fu_7439_p2 = (add_ln703_899_fu_7366_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_834_fu_7444_p2 = (sub_ln703_813_fu_7370_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_835_fu_7449_p2 = (sub_ln703_814_reg_12735 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_836_fu_7453_p2 = (sub_ln703_815_fu_7374_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_837_fu_7458_p2 = (add_ln703_900_fu_7378_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_838_fu_7463_p2 = (sub_ln703_818_reg_12745 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_839_fu_7467_p2 = (add_ln703_901_fu_7390_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_83_fu_1218_p2 = (sub_ln703_70_reg_10586 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_840_fu_7472_p2 = (add_ln703_902_fu_7394_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_841_fu_7485_p2 = (sub_ln703_822_fu_7398_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_842_fu_7498_p2 = (add_ln703_903_fu_7402_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_843_fu_7503_p2 = (sub_ln703_826_fu_7407_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_844_fu_7508_p2 = (sub_ln703_827_fu_7412_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_845_fu_7518_p2 = (sub_ln703_829_fu_7422_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_846_fu_7523_p2 = (sub_ln703_831_fu_7430_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_847_fu_7528_p2 = (add_ln703_906_reg_12775 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_848_fu_7551_p2 = (sub_ln703_834_fu_7444_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_849_fu_7556_p2 = (sub_ln703_836_fu_7453_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_84_fu_1222_p2 = (add_ln703_177_reg_10591 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_850_fu_7566_p2 = (sub_ln703_839_fu_7467_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_851_fu_7571_p2 = (add_ln703_907_fu_7477_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_852_fu_7319_p2 = (add_ln703_910_fu_7259_p2 - data_57_V_read_3_reg_8786_pp0_iter14_reg);

assign sub_ln703_853_fu_7576_p2 = (add_ln703_911_fu_7481_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_854_fu_7586_p2 = (add_ln703_912_fu_7490_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_855_fu_7591_p2 = (add_ln703_913_fu_7494_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_856_fu_7596_p2 = (add_ln703_917_reg_12780 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_857_fu_7600_p2 = (sub_ln703_842_fu_7498_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_858_fu_7605_p2 = (sub_ln703_843_fu_7503_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_859_fu_7615_p2 = (add_ln703_918_fu_7513_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_85_fu_1230_p2 = (add_ln703_181_reg_10601 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_860_fu_7620_p2 = (sub_ln703_845_fu_7518_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_861_fu_7625_p2 = (add_ln703_922_reg_12785 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_862_fu_7324_p2 = (add_ln703_925_fu_7302_p2 - data_58_V_read_3_reg_8756_pp0_iter14_reg);

assign sub_ln703_863_fu_7639_p2 = (add_ln703_926_fu_7532_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_864_fu_7644_p2 = (add_ln703_928_fu_7541_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_865_fu_7649_p2 = (add_ln703_929_fu_7546_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_866_fu_7654_p2 = (sub_ln703_848_fu_7551_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_867_fu_7669_p2 = (sub_ln703_849_fu_7556_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_868_fu_7674_p2 = (add_ln703_930_fu_7561_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_869_fu_7329_p2 = (add_ln703_932_fu_7313_p2 - data_58_V_read_3_reg_8756_pp0_iter14_reg);

assign sub_ln703_86_fu_1234_p2 = (add_ln703_183_reg_10606 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_870_fu_7685_p2 = (sub_ln703_850_fu_7566_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_871_fu_7696_p2 = (sub_ln703_851_fu_7571_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_872_fu_7705_p2 = (sub_ln703_853_fu_7576_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_873_fu_7710_p2 = (add_ln703_933_fu_7581_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_874_fu_7725_p2 = (sub_ln703_855_fu_7591_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_875_fu_7730_p2 = (sub_ln703_856_fu_7596_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_876_fu_7878_p2 = (sub_ln703_857_reg_12835 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_877_fu_7886_p2 = (add_ln703_934_reg_12845 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_878_fu_7890_p2 = (sub_ln703_859_reg_12850 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_879_fu_7735_p2 = (sub_ln703_860_fu_7620_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_87_fu_1238_p2 = (add_ln703_184_fu_1143_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_880_fu_7750_p2 = (sub_ln703_861_fu_7625_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_881_fu_7755_p2 = (add_ln703_935_fu_7629_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_882_fu_7894_p2 = (add_ln703_936_reg_12855 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_883_fu_7898_p2 = (sub_ln703_863_reg_12860 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_884_fu_7902_p2 = (sub_ln703_865_reg_12865 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_885_fu_7906_p2 = (sub_ln703_866_reg_12870 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_886_fu_7910_p2 = (add_ln703_938_reg_12875 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_887_fu_7914_p2 = (sub_ln703_867_reg_12880 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_888_fu_7918_p2 = (sub_ln703_868_reg_12885 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_889_fu_7922_p2 = (sub_ln703_869_reg_12800_pp0_iter16_reg - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_88_fu_1248_p2 = (sub_ln703_73_reg_10611 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_890_fu_7926_p2 = (add_ln703_939_reg_12890 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_891_fu_7930_p2 = (sub_ln703_870_reg_12895 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_892_fu_7780_p2 = (add_ln703_940_fu_7690_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_893_fu_7785_p2 = (sub_ln703_871_fu_7696_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_894_fu_7790_p2 = (add_ln703_941_fu_7701_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_895_fu_7795_p2 = (sub_ln703_872_fu_7705_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_896_fu_7934_p2 = (sub_ln703_873_reg_12900 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_897_fu_7938_p2 = (add_ln703_943_reg_12905 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_898_fu_7805_p2 = (sub_ln703_874_fu_7725_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_899_fu_7942_p2 = (sub_ln703_875_reg_12910 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_89_fu_1252_p2 = (sub_ln703_74_fu_1151_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_8_fu_572_p2 = (sub_ln703_4_reg_10361 - data_3_V_read_10_reg_10295_pp0_iter1_reg);

assign sub_ln703_900_fu_7946_p2 = (sub_ln703_876_fu_7878_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_901_fu_7951_p2 = (add_ln703_944_fu_7882_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_902_fu_7961_p2 = (sub_ln703_878_fu_7890_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_903_fu_7966_p2 = (sub_ln703_879_reg_12915 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_904_fu_7810_p2 = (add_ln703_947_fu_7745_p2 - data_60_V_read61_reg_8691_pp0_iter15_reg);

assign sub_ln703_905_fu_7970_p2 = (sub_ln703_880_reg_12920 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_906_fu_7974_p2 = (sub_ln703_881_reg_12925 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_907_fu_7978_p2 = (sub_ln703_883_fu_7898_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_908_fu_7983_p2 = (add_ln703_948_reg_12930 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_909_fu_7987_p2 = (sub_ln703_885_fu_7906_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_90_fu_1257_p2 = (sub_ln703_75_reg_10616 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_910_fu_7992_p2 = (sub_ln703_888_fu_7918_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_911_fu_7833_p2 = (add_ln703_951_fu_7774_p2 - data_60_V_read61_reg_8691_pp0_iter15_reg);

assign sub_ln703_912_fu_8002_p2 = (sub_ln703_890_fu_7926_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_913_fu_8007_p2 = (sub_ln703_891_fu_7930_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_914_fu_8020_p2 = (sub_ln703_894_reg_12945 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_915_fu_8024_p2 = (sub_ln703_895_reg_12950 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_916_fu_8028_p2 = (sub_ln703_896_fu_7934_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_917_fu_7838_p2 = (add_ln703_952_fu_7800_p2 - data_60_V_read61_reg_8691_pp0_iter15_reg);

assign sub_ln703_918_fu_8033_p2 = (sub_ln703_898_reg_12955 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_919_fu_8037_p2 = (add_ln703_953_fu_7956_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_91_fu_1261_p2 = (add_ln703_186_reg_10621 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_920_fu_8042_p2 = (sub_ln703_902_fu_7961_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_921_fu_8047_p2 = (sub_ln703_903_fu_7966_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_922_fu_7843_p2 = (add_ln703_955_fu_7815_p2 - data_61_V_read62_reg_8663_pp0_iter15_reg);

assign sub_ln703_923_fu_8057_p2 = (sub_ln703_906_fu_7974_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_924_fu_8072_p2 = (add_ln703_958_reg_12965 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_925_fu_8076_p2 = (sub_ln703_911_reg_12970 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_926_fu_8080_p2 = (add_ln703_959_fu_7997_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_927_fu_8085_p2 = (sub_ln703_913_fu_8007_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_928_fu_8090_p2 = (add_ln703_960_fu_8012_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_929_fu_8095_p2 = (add_ln703_961_fu_8016_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_92_fu_1054_p2 = (add_ln703_189_fu_1045_p2 - data_9_V_read_8_reg_10136_pp0_iter3_reg);

assign sub_ln703_930_fu_8120_p2 = (sub_ln703_921_fu_8047_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_931_fu_8134_p2 = (add_ln703_962_fu_8052_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_932_fu_8139_p2 = (sub_ln703_922_reg_12980 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_933_fu_8143_p2 = (sub_ln703_923_fu_8057_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_934_fu_8165_p2 = (add_ln703_963_fu_8062_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_935_fu_8181_p2 = (add_ln703_965_fu_8067_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_936_fu_8209_p2 = (sub_ln703_928_fu_8090_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_937_fu_8219_p2 = (add_ln703_966_fu_8100_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_938_fu_8224_p2 = (add_ln703_967_fu_8105_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_939_fu_8229_p2 = (add_ln703_968_fu_8110_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_93_fu_1275_p2 = (sub_ln703_79_fu_1168_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_940_fu_8234_p2 = (add_ln703_969_fu_8115_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_94_fu_1280_p2 = (add_ln703_190_fu_1172_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_95_fu_1285_p2 = (add_ln703_191_fu_1176_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_96_fu_1294_p2 = (add_ln703_193_fu_1180_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_97_fu_1304_p2 = (add_ln703_194_fu_1189_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_98_fu_1319_p2 = (add_ln703_195_fu_1204_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_99_fu_1324_p2 = (add_ln703_197_fu_1209_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_9_fu_611_p2 = (sub_ln703_3_reg_10379 - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_fu_536_p2 = (data_1_V_read_10_reg_10323 - data_0_V_read_10_reg_10329);

endmodule //dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;

reg   [15:0] data_31_V_read32_reg_989;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter1_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter2_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter3_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter4_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter5_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter6_reg;
reg   [15:0] data_30_V_read31_reg_998;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter1_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter2_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter3_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter4_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter5_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter6_reg;
reg   [15:0] data_29_V_read_6_reg_1006;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter1_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter2_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter3_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter4_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter5_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter6_reg;
reg   [15:0] data_28_V_read_6_reg_1014;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter1_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter2_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter3_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter4_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter5_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter6_reg;
reg   [15:0] data_27_V_read_7_reg_1023;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter1_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter2_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter3_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter4_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter5_reg;
reg   [15:0] data_26_V_read_7_reg_1032;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter1_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter2_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter3_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter4_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter5_reg;
reg   [15:0] data_25_V_read26_reg_1041;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter1_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter2_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter3_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter4_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter5_reg;
reg   [15:0] data_24_V_read25_reg_1050;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter1_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter2_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter3_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter4_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter5_reg;
reg   [15:0] data_23_V_read24_reg_1059;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter1_reg;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter2_reg;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter3_reg;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_1068;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter1_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter2_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter3_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter5_reg;
reg   [15:0] data_21_V_read22_reg_1077;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter1_reg;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter2_reg;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter3_reg;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter4_reg;
reg   [15:0] data_20_V_read21_reg_1086;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter1_reg;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter2_reg;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter3_reg;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter4_reg;
reg   [15:0] data_19_V_read_6_reg_1095;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter1_reg;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter2_reg;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter3_reg;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter4_reg;
reg   [15:0] data_18_V_read_6_reg_1103;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter1_reg;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter2_reg;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter3_reg;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter4_reg;
reg   [15:0] data_17_V_read_7_reg_1111;
reg   [15:0] data_17_V_read_7_reg_1111_pp0_iter1_reg;
reg   [15:0] data_17_V_read_7_reg_1111_pp0_iter2_reg;
reg   [15:0] data_17_V_read_7_reg_1111_pp0_iter3_reg;
reg   [15:0] data_16_V_read_7_reg_1120;
reg   [15:0] data_16_V_read_7_reg_1120_pp0_iter1_reg;
reg   [15:0] data_16_V_read_7_reg_1120_pp0_iter2_reg;
reg   [15:0] data_16_V_read_7_reg_1120_pp0_iter3_reg;
reg   [15:0] data_15_V_read16_reg_1129;
reg   [15:0] data_15_V_read16_reg_1129_pp0_iter1_reg;
reg   [15:0] data_15_V_read16_reg_1129_pp0_iter2_reg;
reg   [15:0] data_15_V_read16_reg_1129_pp0_iter3_reg;
reg   [15:0] data_14_V_read15_reg_1138;
reg   [15:0] data_14_V_read15_reg_1138_pp0_iter1_reg;
reg   [15:0] data_14_V_read15_reg_1138_pp0_iter2_reg;
reg   [15:0] data_14_V_read15_reg_1138_pp0_iter3_reg;
reg   [15:0] data_13_V_read14_reg_1147;
reg   [15:0] data_13_V_read14_reg_1147_pp0_iter1_reg;
reg   [15:0] data_13_V_read14_reg_1147_pp0_iter2_reg;
reg   [15:0] data_12_V_read13_reg_1156;
reg   [15:0] data_12_V_read13_reg_1156_pp0_iter1_reg;
reg   [15:0] data_12_V_read13_reg_1156_pp0_iter2_reg;
reg   [15:0] data_11_V_read12_reg_1165;
reg   [15:0] data_11_V_read12_reg_1165_pp0_iter1_reg;
reg   [15:0] data_11_V_read12_reg_1165_pp0_iter2_reg;
reg   [15:0] data_10_V_read11_reg_1174;
reg   [15:0] data_10_V_read11_reg_1174_pp0_iter1_reg;
reg   [15:0] data_10_V_read11_reg_1174_pp0_iter2_reg;
reg   [15:0] data_9_V_read_6_reg_1183;
reg   [15:0] data_9_V_read_6_reg_1183_pp0_iter1_reg;
reg   [15:0] data_8_V_read_6_reg_1192;
reg   [15:0] data_8_V_read_6_reg_1192_pp0_iter1_reg;
reg   [15:0] data_7_V_read_7_reg_1201;
reg   [15:0] data_7_V_read_7_reg_1201_pp0_iter1_reg;
reg   [15:0] data_6_V_read_7_reg_1208;
reg   [15:0] data_5_V_read_7_reg_1215;
reg   [15:0] data_5_V_read_7_reg_1215_pp0_iter1_reg;
reg   [15:0] data_4_V_read_8_reg_1224;
reg   [15:0] data_3_V_read_8_reg_1232;
reg   [15:0] data_2_V_read_8_reg_1240;
wire   [15:0] add_ln703_fu_280_p2;
reg   [15:0] add_ln703_reg_1246;
wire   [15:0] sub_ln703_1_fu_286_p2;
reg   [15:0] sub_ln703_1_reg_1252;
wire   [15:0] sub_ln703_5_fu_319_p2;
reg   [15:0] sub_ln703_5_reg_1258;
wire   [15:0] sub_ln703_6_fu_324_p2;
reg   [15:0] sub_ln703_6_reg_1263;
wire   [15:0] add_ln703_136_fu_347_p2;
reg   [15:0] add_ln703_136_reg_1268;
wire   [15:0] sub_ln703_9_fu_353_p2;
reg   [15:0] sub_ln703_9_reg_1273;
wire   [15:0] add_ln703_138_fu_363_p2;
reg   [15:0] add_ln703_138_reg_1278;
wire   [15:0] add_ln703_139_fu_367_p2;
reg   [15:0] add_ln703_139_reg_1284;
wire   [15:0] add_ln703_145_fu_433_p2;
reg   [15:0] add_ln703_145_reg_1289;
wire   [15:0] sub_ln703_18_fu_443_p2;
reg   [15:0] sub_ln703_18_reg_1294;
wire   [15:0] add_ln703_146_fu_453_p2;
reg   [15:0] add_ln703_146_reg_1299;
wire   [15:0] add_ln703_147_fu_458_p2;
reg   [15:0] add_ln703_147_reg_1304;
wire   [15:0] add_ln703_148_fu_463_p2;
reg   [15:0] add_ln703_148_reg_1309;
wire   [15:0] add_ln703_149_fu_468_p2;
reg   [15:0] add_ln703_149_reg_1314;
wire   [15:0] sub_ln703_25_fu_517_p2;
reg   [15:0] sub_ln703_25_reg_1319;
wire   [15:0] sub_ln703_26_fu_527_p2;
reg   [15:0] sub_ln703_26_reg_1324;
wire   [15:0] sub_ln703_28_fu_537_p2;
reg   [15:0] sub_ln703_28_reg_1329;
wire   [15:0] sub_ln703_30_fu_542_p2;
reg   [15:0] sub_ln703_30_reg_1334;
wire   [15:0] sub_ln703_33_fu_562_p2;
reg   [15:0] sub_ln703_33_reg_1339;
wire   [15:0] add_ln703_166_fu_567_p2;
reg   [15:0] add_ln703_166_reg_1344;
wire   [15:0] add_ln703_163_fu_621_p2;
reg   [15:0] add_ln703_163_reg_1350;
wire   [15:0] sub_ln703_38_fu_626_p2;
reg   [15:0] sub_ln703_38_reg_1355;
wire   [15:0] add_ln703_167_fu_641_p2;
reg   [15:0] add_ln703_167_reg_1360;
wire   [15:0] sub_ln703_41_fu_646_p2;
reg   [15:0] sub_ln703_41_reg_1365;
wire   [15:0] add_ln703_176_fu_660_p2;
reg   [15:0] add_ln703_176_reg_1370;
reg   [15:0] add_ln703_176_reg_1370_pp0_iter5_reg;
wire   [15:0] sub_ln703_46_fu_697_p2;
reg   [15:0] sub_ln703_46_reg_1375;
wire   [15:0] add_ln703_173_fu_732_p2;
reg   [15:0] add_ln703_173_reg_1380;
wire   [15:0] sub_ln703_49_fu_737_p2;
reg   [15:0] sub_ln703_49_reg_1385;
wire   [15:0] sub_ln703_50_fu_742_p2;
reg   [15:0] sub_ln703_50_reg_1390;
wire   [15:0] add_ln703_180_fu_760_p2;
reg   [15:0] add_ln703_180_reg_1395;
wire   [15:0] add_ln703_184_fu_770_p2;
reg   [15:0] add_ln703_184_reg_1400;
wire   [15:0] sub_ln703_61_fu_840_p2;
reg   [15:0] sub_ln703_61_reg_1405;
wire   [15:0] add_ln703_189_fu_855_p2;
reg   [15:0] add_ln703_189_reg_1410;
wire   [15:0] sub_ln703_62_fu_860_p2;
reg   [15:0] sub_ln703_62_reg_1415;
wire   [15:0] sub_ln703_64_fu_865_p2;
reg   [15:0] sub_ln703_64_reg_1420;
wire   [15:0] add_ln703_192_fu_870_p2;
reg   [15:0] add_ln703_192_reg_1425;
wire   [15:0] add_ln703_194_fu_874_p2;
reg   [15:0] add_ln703_194_reg_1431;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_fu_274_p2;
wire   [15:0] add_ln703_130_fu_300_p2;
wire   [15:0] sub_ln703_2_fu_292_p2;
wire   [15:0] sub_ln703_3_fu_296_p2;
wire   [15:0] add_ln703_131_fu_304_p2;
wire   [15:0] sub_ln703_4_fu_309_p2;
wire   [15:0] add_ln703_132_fu_314_p2;
wire   [15:0] add_ln703_134_fu_338_p2;
wire   [15:0] add_ln703_135_fu_342_p2;
wire   [15:0] add_ln703_133_fu_334_p2;
wire   [15:0] sub_ln703_8_fu_329_p2;
wire   [15:0] add_ln703_137_fu_358_p2;
wire   [15:0] sub_ln703_7_fu_373_p2;
wire   [15:0] add_ln703_141_fu_386_p2;
wire   [15:0] sub_ln703_10_fu_377_p2;
wire   [15:0] add_ln703_140_fu_381_p2;
wire   [15:0] add_ln703_142_fu_390_p2;
wire   [15:0] add_ln703_143_fu_395_p2;
wire   [15:0] add_ln703_144_fu_399_p2;
wire   [15:0] sub_ln703_11_fu_404_p2;
wire   [15:0] sub_ln703_13_fu_413_p2;
wire   [15:0] sub_ln703_14_fu_418_p2;
wire   [15:0] sub_ln703_15_fu_423_p2;
wire   [15:0] sub_ln703_16_fu_428_p2;
wire   [15:0] sub_ln703_17_fu_438_p2;
wire   [15:0] sub_ln703_19_fu_448_p2;
wire   [15:0] sub_ln703_12_fu_408_p2;
wire   [15:0] sub_ln703_20_fu_472_p2;
wire   [15:0] add_ln703_151_fu_489_p2;
wire   [15:0] add_ln703_150_fu_476_p2;
wire   [15:0] sub_ln703_21_fu_480_p2;
wire   [15:0] sub_ln703_22_fu_485_p2;
wire   [15:0] add_ln703_152_fu_493_p2;
wire   [15:0] sub_ln703_24_fu_502_p2;
wire   [15:0] add_ln703_153_fu_507_p2;
wire   [15:0] add_ln703_154_fu_512_p2;
wire   [15:0] add_ln703_155_fu_522_p2;
wire   [15:0] sub_ln703_27_fu_532_p2;
wire   [15:0] sub_ln703_23_fu_498_p2;
wire   [15:0] add_ln703_158_fu_552_p2;
wire   [15:0] add_ln703_157_fu_547_p2;
wire   [15:0] add_ln703_159_fu_556_p2;
wire   [15:0] add_ln703_156_fu_571_p2;
wire   [15:0] sub_ln703_29_fu_575_p2;
wire   [15:0] sub_ln703_32_fu_584_p2;
wire   [15:0] add_ln703_160_fu_588_p2;
wire   [15:0] add_ln703_161_fu_593_p2;
wire   [15:0] sub_ln703_34_fu_597_p2;
wire   [15:0] sub_ln703_35_fu_602_p2;
wire   [15:0] add_ln703_162_fu_616_p2;
wire   [15:0] add_ln703_164_fu_631_p2;
wire   [15:0] sub_ln703_36_fu_607_p2;
wire   [15:0] sub_ln703_37_fu_612_p2;
wire   [15:0] add_ln703_165_fu_635_p2;
wire   [15:0] sub_ln703_31_fu_579_p2;
wire   [15:0] add_ln703_175_fu_656_p2;
wire   [15:0] add_ln703_174_fu_651_p2;
wire   [15:0] sub_ln703_39_fu_666_p2;
wire   [15:0] add_ln703_168_fu_674_p2;
wire   [15:0] sub_ln703_42_fu_679_p2;
wire   [15:0] sub_ln703_43_fu_683_p2;
wire   [15:0] sub_ln703_44_fu_688_p2;
wire   [15:0] sub_ln703_45_fu_692_p2;
wire   [15:0] sub_ln703_40_fu_670_p2;
wire   [15:0] add_ln703_171_fu_717_p2;
wire   [15:0] add_ln703_170_fu_712_p2;
wire   [15:0] add_ln703_169_fu_702_p2;
wire   [15:0] sub_ln703_47_fu_707_p2;
wire   [15:0] add_ln703_172_fu_721_p2;
wire   [15:0] sub_ln703_48_fu_727_p2;
wire   [15:0] add_ln703_178_fu_751_p2;
wire   [15:0] add_ln703_179_fu_755_p2;
wire   [15:0] add_ln703_177_fu_747_p2;
wire   [15:0] add_ln703_183_fu_766_p2;
wire   [15:0] add_ln703_181_fu_775_p2;
wire   [15:0] sub_ln703_51_fu_779_p2;
wire   [15:0] sub_ln703_52_fu_783_p2;
wire   [15:0] add_ln703_182_fu_806_p2;
wire   [15:0] sub_ln703_53_fu_787_p2;
wire   [15:0] sub_ln703_54_fu_791_p2;
wire   [15:0] sub_ln703_56_fu_801_p2;
wire   [15:0] add_ln703_185_fu_810_p2;
wire   [15:0] add_ln703_186_fu_815_p2;
wire   [15:0] sub_ln703_57_fu_820_p2;
wire   [15:0] add_ln703_187_fu_845_p2;
wire   [15:0] sub_ln703_55_fu_796_p2;
wire   [15:0] sub_ln703_59_fu_830_p2;
wire   [15:0] sub_ln703_60_fu_835_p2;
wire   [15:0] add_ln703_188_fu_849_p2;
wire   [15:0] sub_ln703_58_fu_825_p2;
wire   [15:0] sub_ln703_63_fu_879_p2;
wire   [15:0] sub_ln703_65_fu_883_p2;
wire   [15:0] add_ln703_190_fu_887_p2;
wire   [15:0] sub_ln703_66_fu_891_p2;
wire   [15:0] add_ln703_195_fu_915_p2;
wire   [15:0] add_ln703_191_fu_896_p2;
wire   [15:0] sub_ln703_68_fu_906_p2;
wire   [15:0] add_ln703_193_fu_911_p2;
wire   [15:0] add_ln703_196_fu_919_p2;
wire   [15:0] sub_ln703_69_fu_924_p2;
wire   [15:0] add_ln703_198_fu_949_p2;
wire   [15:0] sub_ln703_67_fu_901_p2;
wire   [15:0] sub_ln703_70_fu_929_p2;
wire   [15:0] acc_1_V_fu_934_p2;
wire   [15:0] acc_2_V_fu_939_p2;
wire   [15:0] acc_3_V_fu_944_p2;
wire   [15:0] acc_4_V_fu_953_p2;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln703_136_reg_1268 <= add_ln703_136_fu_347_p2;
        add_ln703_138_reg_1278 <= add_ln703_138_fu_363_p2;
        add_ln703_139_reg_1284 <= add_ln703_139_fu_367_p2;
        add_ln703_145_reg_1289 <= add_ln703_145_fu_433_p2;
        add_ln703_146_reg_1299 <= add_ln703_146_fu_453_p2;
        add_ln703_147_reg_1304 <= add_ln703_147_fu_458_p2;
        add_ln703_148_reg_1309 <= add_ln703_148_fu_463_p2;
        add_ln703_149_reg_1314 <= add_ln703_149_fu_468_p2;
        add_ln703_163_reg_1350 <= add_ln703_163_fu_621_p2;
        add_ln703_166_reg_1344 <= add_ln703_166_fu_567_p2;
        add_ln703_167_reg_1360 <= add_ln703_167_fu_641_p2;
        add_ln703_173_reg_1380 <= add_ln703_173_fu_732_p2;
        add_ln703_176_reg_1370 <= add_ln703_176_fu_660_p2;
        add_ln703_176_reg_1370_pp0_iter5_reg <= add_ln703_176_reg_1370;
        add_ln703_180_reg_1395 <= add_ln703_180_fu_760_p2;
        add_ln703_184_reg_1400 <= add_ln703_184_fu_770_p2;
        add_ln703_189_reg_1410 <= add_ln703_189_fu_855_p2;
        add_ln703_192_reg_1425 <= add_ln703_192_fu_870_p2;
        add_ln703_194_reg_1431 <= add_ln703_194_fu_874_p2;
        add_ln703_reg_1246 <= add_ln703_fu_280_p2;
        data_10_V_read11_reg_1174 <= data_10_V_read_int_reg;
        data_10_V_read11_reg_1174_pp0_iter1_reg <= data_10_V_read11_reg_1174;
        data_10_V_read11_reg_1174_pp0_iter2_reg <= data_10_V_read11_reg_1174_pp0_iter1_reg;
        data_11_V_read12_reg_1165 <= data_11_V_read_int_reg;
        data_11_V_read12_reg_1165_pp0_iter1_reg <= data_11_V_read12_reg_1165;
        data_11_V_read12_reg_1165_pp0_iter2_reg <= data_11_V_read12_reg_1165_pp0_iter1_reg;
        data_12_V_read13_reg_1156 <= data_12_V_read_int_reg;
        data_12_V_read13_reg_1156_pp0_iter1_reg <= data_12_V_read13_reg_1156;
        data_12_V_read13_reg_1156_pp0_iter2_reg <= data_12_V_read13_reg_1156_pp0_iter1_reg;
        data_13_V_read14_reg_1147 <= data_13_V_read_int_reg;
        data_13_V_read14_reg_1147_pp0_iter1_reg <= data_13_V_read14_reg_1147;
        data_13_V_read14_reg_1147_pp0_iter2_reg <= data_13_V_read14_reg_1147_pp0_iter1_reg;
        data_14_V_read15_reg_1138 <= data_14_V_read_int_reg;
        data_14_V_read15_reg_1138_pp0_iter1_reg <= data_14_V_read15_reg_1138;
        data_14_V_read15_reg_1138_pp0_iter2_reg <= data_14_V_read15_reg_1138_pp0_iter1_reg;
        data_14_V_read15_reg_1138_pp0_iter3_reg <= data_14_V_read15_reg_1138_pp0_iter2_reg;
        data_15_V_read16_reg_1129 <= data_15_V_read_int_reg;
        data_15_V_read16_reg_1129_pp0_iter1_reg <= data_15_V_read16_reg_1129;
        data_15_V_read16_reg_1129_pp0_iter2_reg <= data_15_V_read16_reg_1129_pp0_iter1_reg;
        data_15_V_read16_reg_1129_pp0_iter3_reg <= data_15_V_read16_reg_1129_pp0_iter2_reg;
        data_16_V_read_7_reg_1120 <= data_16_V_read_int_reg;
        data_16_V_read_7_reg_1120_pp0_iter1_reg <= data_16_V_read_7_reg_1120;
        data_16_V_read_7_reg_1120_pp0_iter2_reg <= data_16_V_read_7_reg_1120_pp0_iter1_reg;
        data_16_V_read_7_reg_1120_pp0_iter3_reg <= data_16_V_read_7_reg_1120_pp0_iter2_reg;
        data_17_V_read_7_reg_1111 <= data_17_V_read_int_reg;
        data_17_V_read_7_reg_1111_pp0_iter1_reg <= data_17_V_read_7_reg_1111;
        data_17_V_read_7_reg_1111_pp0_iter2_reg <= data_17_V_read_7_reg_1111_pp0_iter1_reg;
        data_17_V_read_7_reg_1111_pp0_iter3_reg <= data_17_V_read_7_reg_1111_pp0_iter2_reg;
        data_18_V_read_6_reg_1103 <= data_18_V_read_int_reg;
        data_18_V_read_6_reg_1103_pp0_iter1_reg <= data_18_V_read_6_reg_1103;
        data_18_V_read_6_reg_1103_pp0_iter2_reg <= data_18_V_read_6_reg_1103_pp0_iter1_reg;
        data_18_V_read_6_reg_1103_pp0_iter3_reg <= data_18_V_read_6_reg_1103_pp0_iter2_reg;
        data_18_V_read_6_reg_1103_pp0_iter4_reg <= data_18_V_read_6_reg_1103_pp0_iter3_reg;
        data_19_V_read_6_reg_1095 <= data_19_V_read_int_reg;
        data_19_V_read_6_reg_1095_pp0_iter1_reg <= data_19_V_read_6_reg_1095;
        data_19_V_read_6_reg_1095_pp0_iter2_reg <= data_19_V_read_6_reg_1095_pp0_iter1_reg;
        data_19_V_read_6_reg_1095_pp0_iter3_reg <= data_19_V_read_6_reg_1095_pp0_iter2_reg;
        data_19_V_read_6_reg_1095_pp0_iter4_reg <= data_19_V_read_6_reg_1095_pp0_iter3_reg;
        data_20_V_read21_reg_1086 <= data_20_V_read_int_reg;
        data_20_V_read21_reg_1086_pp0_iter1_reg <= data_20_V_read21_reg_1086;
        data_20_V_read21_reg_1086_pp0_iter2_reg <= data_20_V_read21_reg_1086_pp0_iter1_reg;
        data_20_V_read21_reg_1086_pp0_iter3_reg <= data_20_V_read21_reg_1086_pp0_iter2_reg;
        data_20_V_read21_reg_1086_pp0_iter4_reg <= data_20_V_read21_reg_1086_pp0_iter3_reg;
        data_21_V_read22_reg_1077 <= data_21_V_read_int_reg;
        data_21_V_read22_reg_1077_pp0_iter1_reg <= data_21_V_read22_reg_1077;
        data_21_V_read22_reg_1077_pp0_iter2_reg <= data_21_V_read22_reg_1077_pp0_iter1_reg;
        data_21_V_read22_reg_1077_pp0_iter3_reg <= data_21_V_read22_reg_1077_pp0_iter2_reg;
        data_21_V_read22_reg_1077_pp0_iter4_reg <= data_21_V_read22_reg_1077_pp0_iter3_reg;
        data_22_V_read23_reg_1068 <= data_22_V_read_int_reg;
        data_22_V_read23_reg_1068_pp0_iter1_reg <= data_22_V_read23_reg_1068;
        data_22_V_read23_reg_1068_pp0_iter2_reg <= data_22_V_read23_reg_1068_pp0_iter1_reg;
        data_22_V_read23_reg_1068_pp0_iter3_reg <= data_22_V_read23_reg_1068_pp0_iter2_reg;
        data_22_V_read23_reg_1068_pp0_iter4_reg <= data_22_V_read23_reg_1068_pp0_iter3_reg;
        data_22_V_read23_reg_1068_pp0_iter5_reg <= data_22_V_read23_reg_1068_pp0_iter4_reg;
        data_23_V_read24_reg_1059 <= data_23_V_read_int_reg;
        data_23_V_read24_reg_1059_pp0_iter1_reg <= data_23_V_read24_reg_1059;
        data_23_V_read24_reg_1059_pp0_iter2_reg <= data_23_V_read24_reg_1059_pp0_iter1_reg;
        data_23_V_read24_reg_1059_pp0_iter3_reg <= data_23_V_read24_reg_1059_pp0_iter2_reg;
        data_23_V_read24_reg_1059_pp0_iter4_reg <= data_23_V_read24_reg_1059_pp0_iter3_reg;
        data_24_V_read25_reg_1050 <= data_24_V_read_int_reg;
        data_24_V_read25_reg_1050_pp0_iter1_reg <= data_24_V_read25_reg_1050;
        data_24_V_read25_reg_1050_pp0_iter2_reg <= data_24_V_read25_reg_1050_pp0_iter1_reg;
        data_24_V_read25_reg_1050_pp0_iter3_reg <= data_24_V_read25_reg_1050_pp0_iter2_reg;
        data_24_V_read25_reg_1050_pp0_iter4_reg <= data_24_V_read25_reg_1050_pp0_iter3_reg;
        data_24_V_read25_reg_1050_pp0_iter5_reg <= data_24_V_read25_reg_1050_pp0_iter4_reg;
        data_25_V_read26_reg_1041 <= data_25_V_read_int_reg;
        data_25_V_read26_reg_1041_pp0_iter1_reg <= data_25_V_read26_reg_1041;
        data_25_V_read26_reg_1041_pp0_iter2_reg <= data_25_V_read26_reg_1041_pp0_iter1_reg;
        data_25_V_read26_reg_1041_pp0_iter3_reg <= data_25_V_read26_reg_1041_pp0_iter2_reg;
        data_25_V_read26_reg_1041_pp0_iter4_reg <= data_25_V_read26_reg_1041_pp0_iter3_reg;
        data_25_V_read26_reg_1041_pp0_iter5_reg <= data_25_V_read26_reg_1041_pp0_iter4_reg;
        data_26_V_read_7_reg_1032 <= data_26_V_read_int_reg;
        data_26_V_read_7_reg_1032_pp0_iter1_reg <= data_26_V_read_7_reg_1032;
        data_26_V_read_7_reg_1032_pp0_iter2_reg <= data_26_V_read_7_reg_1032_pp0_iter1_reg;
        data_26_V_read_7_reg_1032_pp0_iter3_reg <= data_26_V_read_7_reg_1032_pp0_iter2_reg;
        data_26_V_read_7_reg_1032_pp0_iter4_reg <= data_26_V_read_7_reg_1032_pp0_iter3_reg;
        data_26_V_read_7_reg_1032_pp0_iter5_reg <= data_26_V_read_7_reg_1032_pp0_iter4_reg;
        data_27_V_read_7_reg_1023 <= data_27_V_read_int_reg;
        data_27_V_read_7_reg_1023_pp0_iter1_reg <= data_27_V_read_7_reg_1023;
        data_27_V_read_7_reg_1023_pp0_iter2_reg <= data_27_V_read_7_reg_1023_pp0_iter1_reg;
        data_27_V_read_7_reg_1023_pp0_iter3_reg <= data_27_V_read_7_reg_1023_pp0_iter2_reg;
        data_27_V_read_7_reg_1023_pp0_iter4_reg <= data_27_V_read_7_reg_1023_pp0_iter3_reg;
        data_27_V_read_7_reg_1023_pp0_iter5_reg <= data_27_V_read_7_reg_1023_pp0_iter4_reg;
        data_28_V_read_6_reg_1014 <= data_28_V_read_int_reg;
        data_28_V_read_6_reg_1014_pp0_iter1_reg <= data_28_V_read_6_reg_1014;
        data_28_V_read_6_reg_1014_pp0_iter2_reg <= data_28_V_read_6_reg_1014_pp0_iter1_reg;
        data_28_V_read_6_reg_1014_pp0_iter3_reg <= data_28_V_read_6_reg_1014_pp0_iter2_reg;
        data_28_V_read_6_reg_1014_pp0_iter4_reg <= data_28_V_read_6_reg_1014_pp0_iter3_reg;
        data_28_V_read_6_reg_1014_pp0_iter5_reg <= data_28_V_read_6_reg_1014_pp0_iter4_reg;
        data_28_V_read_6_reg_1014_pp0_iter6_reg <= data_28_V_read_6_reg_1014_pp0_iter5_reg;
        data_29_V_read_6_reg_1006 <= data_29_V_read_int_reg;
        data_29_V_read_6_reg_1006_pp0_iter1_reg <= data_29_V_read_6_reg_1006;
        data_29_V_read_6_reg_1006_pp0_iter2_reg <= data_29_V_read_6_reg_1006_pp0_iter1_reg;
        data_29_V_read_6_reg_1006_pp0_iter3_reg <= data_29_V_read_6_reg_1006_pp0_iter2_reg;
        data_29_V_read_6_reg_1006_pp0_iter4_reg <= data_29_V_read_6_reg_1006_pp0_iter3_reg;
        data_29_V_read_6_reg_1006_pp0_iter5_reg <= data_29_V_read_6_reg_1006_pp0_iter4_reg;
        data_29_V_read_6_reg_1006_pp0_iter6_reg <= data_29_V_read_6_reg_1006_pp0_iter5_reg;
        data_2_V_read_8_reg_1240 <= data_2_V_read_int_reg;
        data_30_V_read31_reg_998 <= data_30_V_read_int_reg;
        data_30_V_read31_reg_998_pp0_iter1_reg <= data_30_V_read31_reg_998;
        data_30_V_read31_reg_998_pp0_iter2_reg <= data_30_V_read31_reg_998_pp0_iter1_reg;
        data_30_V_read31_reg_998_pp0_iter3_reg <= data_30_V_read31_reg_998_pp0_iter2_reg;
        data_30_V_read31_reg_998_pp0_iter4_reg <= data_30_V_read31_reg_998_pp0_iter3_reg;
        data_30_V_read31_reg_998_pp0_iter5_reg <= data_30_V_read31_reg_998_pp0_iter4_reg;
        data_30_V_read31_reg_998_pp0_iter6_reg <= data_30_V_read31_reg_998_pp0_iter5_reg;
        data_31_V_read32_reg_989 <= data_31_V_read_int_reg;
        data_31_V_read32_reg_989_pp0_iter1_reg <= data_31_V_read32_reg_989;
        data_31_V_read32_reg_989_pp0_iter2_reg <= data_31_V_read32_reg_989_pp0_iter1_reg;
        data_31_V_read32_reg_989_pp0_iter3_reg <= data_31_V_read32_reg_989_pp0_iter2_reg;
        data_31_V_read32_reg_989_pp0_iter4_reg <= data_31_V_read32_reg_989_pp0_iter3_reg;
        data_31_V_read32_reg_989_pp0_iter5_reg <= data_31_V_read32_reg_989_pp0_iter4_reg;
        data_31_V_read32_reg_989_pp0_iter6_reg <= data_31_V_read32_reg_989_pp0_iter5_reg;
        data_3_V_read_8_reg_1232 <= data_3_V_read_int_reg;
        data_4_V_read_8_reg_1224 <= data_4_V_read_int_reg;
        data_5_V_read_7_reg_1215 <= data_5_V_read_int_reg;
        data_5_V_read_7_reg_1215_pp0_iter1_reg <= data_5_V_read_7_reg_1215;
        data_6_V_read_7_reg_1208 <= data_6_V_read_int_reg;
        data_7_V_read_7_reg_1201 <= data_7_V_read_int_reg;
        data_7_V_read_7_reg_1201_pp0_iter1_reg <= data_7_V_read_7_reg_1201;
        data_8_V_read_6_reg_1192 <= data_8_V_read_int_reg;
        data_8_V_read_6_reg_1192_pp0_iter1_reg <= data_8_V_read_6_reg_1192;
        data_9_V_read_6_reg_1183 <= data_9_V_read_int_reg;
        data_9_V_read_6_reg_1183_pp0_iter1_reg <= data_9_V_read_6_reg_1183;
        sub_ln703_18_reg_1294 <= sub_ln703_18_fu_443_p2;
        sub_ln703_1_reg_1252 <= sub_ln703_1_fu_286_p2;
        sub_ln703_25_reg_1319 <= sub_ln703_25_fu_517_p2;
        sub_ln703_26_reg_1324 <= sub_ln703_26_fu_527_p2;
        sub_ln703_28_reg_1329 <= sub_ln703_28_fu_537_p2;
        sub_ln703_30_reg_1334 <= sub_ln703_30_fu_542_p2;
        sub_ln703_33_reg_1339 <= sub_ln703_33_fu_562_p2;
        sub_ln703_38_reg_1355 <= sub_ln703_38_fu_626_p2;
        sub_ln703_41_reg_1365 <= sub_ln703_41_fu_646_p2;
        sub_ln703_46_reg_1375 <= sub_ln703_46_fu_697_p2;
        sub_ln703_49_reg_1385 <= sub_ln703_49_fu_737_p2;
        sub_ln703_50_reg_1390 <= sub_ln703_50_fu_742_p2;
        sub_ln703_5_reg_1258 <= sub_ln703_5_fu_319_p2;
        sub_ln703_61_reg_1405 <= sub_ln703_61_fu_840_p2;
        sub_ln703_62_reg_1415 <= sub_ln703_62_fu_860_p2;
        sub_ln703_64_reg_1420 <= sub_ln703_64_fu_865_p2;
        sub_ln703_6_reg_1263 <= sub_ln703_6_fu_324_p2;
        sub_ln703_9_reg_1273 <= sub_ln703_9_fu_353_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= sub_ln703_70_fu_929_p2;
        ap_return_1_int_reg <= acc_1_V_fu_934_p2;
        ap_return_2_int_reg <= acc_2_V_fu_939_p2;
        ap_return_3_int_reg <= acc_3_V_fu_944_p2;
        ap_return_4_int_reg <= acc_4_V_fu_953_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = sub_ln703_70_fu_929_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_934_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_939_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_944_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_953_p2;
    end
end

assign acc_1_V_fu_934_p2 = (add_ln703_193_fu_911_p2 - data_31_V_read32_reg_989_pp0_iter6_reg);

assign acc_2_V_fu_939_p2 = (add_ln703_196_fu_919_p2 - data_31_V_read32_reg_989_pp0_iter6_reg);

assign acc_3_V_fu_944_p2 = (sub_ln703_69_fu_924_p2 + data_31_V_read32_reg_989_pp0_iter6_reg);

assign acc_4_V_fu_953_p2 = (add_ln703_198_fu_949_p2 + sub_ln703_67_fu_901_p2);

assign add_ln703_130_fu_300_p2 = (data_2_V_read_8_reg_1240 + data_3_V_read_8_reg_1232);

assign add_ln703_131_fu_304_p2 = (add_ln703_130_fu_300_p2 + add_ln703_reg_1246);

assign add_ln703_132_fu_314_p2 = (sub_ln703_3_fu_296_p2 + data_4_V_read_8_reg_1224);

assign add_ln703_133_fu_334_p2 = (sub_ln703_1_reg_1252 + data_3_V_read_8_reg_1232);

assign add_ln703_134_fu_338_p2 = (data_5_V_read_7_reg_1215 + data_6_V_read_7_reg_1208);

assign add_ln703_135_fu_342_p2 = (add_ln703_134_fu_338_p2 + data_4_V_read_8_reg_1224);

assign add_ln703_136_fu_347_p2 = (add_ln703_135_fu_342_p2 + add_ln703_133_fu_334_p2);

assign add_ln703_137_fu_358_p2 = (add_ln703_132_fu_314_p2 + data_5_V_read_7_reg_1215);

assign add_ln703_138_fu_363_p2 = (data_6_V_read_7_reg_1208 + data_7_V_read_7_reg_1201);

assign add_ln703_139_fu_367_p2 = (add_ln703_138_fu_363_p2 + add_ln703_137_fu_358_p2);

assign add_ln703_140_fu_381_p2 = (add_ln703_138_reg_1278 + sub_ln703_7_fu_373_p2);

assign add_ln703_141_fu_386_p2 = (sub_ln703_6_reg_1263 + data_5_V_read_7_reg_1215_pp0_iter1_reg);

assign add_ln703_142_fu_390_p2 = (add_ln703_138_reg_1278 + add_ln703_141_fu_386_p2);

assign add_ln703_143_fu_395_p2 = (sub_ln703_9_reg_1273 + data_7_V_read_7_reg_1201_pp0_iter1_reg);

assign add_ln703_144_fu_399_p2 = (sub_ln703_10_fu_377_p2 + data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign add_ln703_145_fu_433_p2 = (sub_ln703_13_fu_413_p2 + data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign add_ln703_146_fu_453_p2 = (sub_ln703_17_fu_438_p2 + data_10_V_read11_reg_1174_pp0_iter1_reg);

assign add_ln703_147_fu_458_p2 = (sub_ln703_19_fu_448_p2 + data_11_V_read12_reg_1165_pp0_iter1_reg);

assign add_ln703_148_fu_463_p2 = (sub_ln703_12_fu_408_p2 + data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign add_ln703_149_fu_468_p2 = (data_10_V_read11_reg_1174_pp0_iter1_reg + data_11_V_read12_reg_1165_pp0_iter1_reg);

assign add_ln703_150_fu_476_p2 = (add_ln703_149_reg_1314 + add_ln703_148_reg_1309);

assign add_ln703_151_fu_489_p2 = (data_11_V_read12_reg_1165_pp0_iter2_reg + data_12_V_read13_reg_1156_pp0_iter2_reg);

assign add_ln703_152_fu_493_p2 = (add_ln703_151_fu_489_p2 + sub_ln703_18_reg_1294);

assign add_ln703_153_fu_507_p2 = (sub_ln703_21_fu_480_p2 + data_12_V_read13_reg_1156_pp0_iter2_reg);

assign add_ln703_154_fu_512_p2 = (sub_ln703_22_fu_485_p2 + data_12_V_read13_reg_1156_pp0_iter2_reg);

assign add_ln703_155_fu_522_p2 = (sub_ln703_24_fu_502_p2 + data_13_V_read14_reg_1147_pp0_iter2_reg);

assign add_ln703_156_fu_571_p2 = (sub_ln703_25_reg_1319 + data_14_V_read15_reg_1138_pp0_iter3_reg);

assign add_ln703_157_fu_547_p2 = (sub_ln703_23_fu_498_p2 + data_13_V_read14_reg_1147_pp0_iter2_reg);

assign add_ln703_158_fu_552_p2 = (data_14_V_read15_reg_1138_pp0_iter2_reg + data_15_V_read16_reg_1129_pp0_iter2_reg);

assign add_ln703_159_fu_556_p2 = (add_ln703_158_fu_552_p2 + add_ln703_157_fu_547_p2);

assign add_ln703_160_fu_588_p2 = (sub_ln703_29_fu_575_p2 + data_15_V_read16_reg_1129_pp0_iter3_reg);

assign add_ln703_161_fu_593_p2 = (sub_ln703_30_reg_1334 + data_15_V_read16_reg_1129_pp0_iter3_reg);

assign add_ln703_162_fu_616_p2 = (sub_ln703_34_fu_597_p2 + data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign add_ln703_163_fu_621_p2 = (sub_ln703_35_fu_602_p2 + data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign add_ln703_164_fu_631_p2 = (data_17_V_read_7_reg_1111_pp0_iter3_reg + data_18_V_read_6_reg_1103_pp0_iter3_reg);

assign add_ln703_165_fu_635_p2 = (add_ln703_164_fu_631_p2 + sub_ln703_36_fu_607_p2);

assign add_ln703_166_fu_567_p2 = (data_18_V_read_6_reg_1103_pp0_iter2_reg + data_19_V_read_6_reg_1095_pp0_iter2_reg);

assign add_ln703_167_fu_641_p2 = (add_ln703_166_reg_1344 + sub_ln703_37_fu_612_p2);

assign add_ln703_168_fu_674_p2 = (sub_ln703_39_fu_666_p2 + data_19_V_read_6_reg_1095_pp0_iter4_reg);

assign add_ln703_169_fu_702_p2 = (sub_ln703_44_fu_688_p2 + data_21_V_read22_reg_1077_pp0_iter4_reg);

assign add_ln703_170_fu_712_p2 = (sub_ln703_40_fu_670_p2 + data_20_V_read21_reg_1086_pp0_iter4_reg);

assign add_ln703_171_fu_717_p2 = (data_21_V_read22_reg_1077_pp0_iter4_reg + data_22_V_read23_reg_1068_pp0_iter4_reg);

assign add_ln703_172_fu_721_p2 = (add_ln703_171_fu_717_p2 + add_ln703_170_fu_712_p2);

assign add_ln703_173_fu_732_p2 = (sub_ln703_47_fu_707_p2 + data_23_V_read24_reg_1059_pp0_iter4_reg);

assign add_ln703_174_fu_651_p2 = (sub_ln703_31_fu_579_p2 + data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign add_ln703_175_fu_656_p2 = (add_ln703_166_reg_1344 + data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign add_ln703_176_fu_660_p2 = (add_ln703_175_fu_656_p2 + add_ln703_174_fu_651_p2);

assign add_ln703_177_fu_747_p2 = (data_20_V_read21_reg_1086_pp0_iter4_reg + data_21_V_read22_reg_1077_pp0_iter4_reg);

assign add_ln703_178_fu_751_p2 = (data_23_V_read24_reg_1059_pp0_iter4_reg + data_24_V_read25_reg_1050_pp0_iter4_reg);

assign add_ln703_179_fu_755_p2 = (add_ln703_178_fu_751_p2 + data_22_V_read23_reg_1068_pp0_iter4_reg);

assign add_ln703_180_fu_760_p2 = (add_ln703_179_fu_755_p2 + add_ln703_177_fu_747_p2);

assign add_ln703_181_fu_775_p2 = (add_ln703_180_reg_1395 + add_ln703_176_reg_1370_pp0_iter5_reg);

assign add_ln703_182_fu_806_p2 = (sub_ln703_46_reg_1375 + data_22_V_read23_reg_1068_pp0_iter5_reg);

assign add_ln703_183_fu_766_p2 = (data_24_V_read25_reg_1050_pp0_iter4_reg + data_25_V_read26_reg_1041_pp0_iter4_reg);

assign add_ln703_184_fu_770_p2 = (add_ln703_183_fu_766_p2 + data_23_V_read24_reg_1059_pp0_iter4_reg);

assign add_ln703_185_fu_810_p2 = (add_ln703_184_reg_1400 + add_ln703_182_fu_806_p2);

assign add_ln703_186_fu_815_p2 = (sub_ln703_53_fu_787_p2 + data_25_V_read26_reg_1041_pp0_iter5_reg);

assign add_ln703_187_fu_845_p2 = (data_26_V_read_7_reg_1032_pp0_iter5_reg + data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign add_ln703_188_fu_849_p2 = (add_ln703_187_fu_845_p2 + sub_ln703_55_fu_796_p2);

assign add_ln703_189_fu_855_p2 = (sub_ln703_59_fu_830_p2 + data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign add_ln703_190_fu_887_p2 = (sub_ln703_62_reg_1415 + data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign add_ln703_191_fu_896_p2 = (sub_ln703_65_fu_883_p2 + data_29_V_read_6_reg_1006_pp0_iter6_reg);

assign add_ln703_192_fu_870_p2 = (data_29_V_read_6_reg_1006_pp0_iter5_reg + data_30_V_read31_reg_998_pp0_iter5_reg);

assign add_ln703_193_fu_911_p2 = (add_ln703_192_reg_1425 + sub_ln703_64_reg_1420);

assign add_ln703_194_fu_874_p2 = (sub_ln703_58_fu_825_p2 + data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign add_ln703_195_fu_915_p2 = (add_ln703_192_reg_1425 + data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign add_ln703_196_fu_919_p2 = (add_ln703_195_fu_915_p2 + add_ln703_194_reg_1431);

assign add_ln703_198_fu_949_p2 = (data_30_V_read31_reg_998_pp0_iter6_reg + data_31_V_read32_reg_989_pp0_iter6_reg);

assign add_ln703_fu_280_p2 = (data_0_V_read_int_reg + data_1_V_read_int_reg);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign sub_ln703_10_fu_377_p2 = (add_ln703_136_reg_1268 - data_7_V_read_7_reg_1201_pp0_iter1_reg);

assign sub_ln703_11_fu_404_p2 = (add_ln703_139_reg_1284 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_12_fu_408_p2 = (add_ln703_140_fu_381_p2 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_13_fu_413_p2 = (add_ln703_142_fu_390_p2 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_14_fu_418_p2 = (add_ln703_143_fu_395_p2 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_15_fu_423_p2 = (add_ln703_144_fu_399_p2 - data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign sub_ln703_16_fu_428_p2 = (sub_ln703_11_fu_404_p2 - data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign sub_ln703_17_fu_438_p2 = (sub_ln703_14_fu_418_p2 - data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign sub_ln703_18_fu_443_p2 = (sub_ln703_15_fu_423_p2 - data_10_V_read11_reg_1174_pp0_iter1_reg);

assign sub_ln703_19_fu_448_p2 = (sub_ln703_16_fu_428_p2 - data_10_V_read11_reg_1174_pp0_iter1_reg);

assign sub_ln703_1_fu_286_p2 = (sub_ln703_fu_274_p2 - data_2_V_read_int_reg);

assign sub_ln703_20_fu_472_p2 = (add_ln703_145_reg_1289 - data_10_V_read11_reg_1174_pp0_iter2_reg);

assign sub_ln703_21_fu_480_p2 = (sub_ln703_20_fu_472_p2 - data_11_V_read12_reg_1165_pp0_iter2_reg);

assign sub_ln703_22_fu_485_p2 = (add_ln703_146_reg_1299 - data_11_V_read12_reg_1165_pp0_iter2_reg);

assign sub_ln703_23_fu_498_p2 = (add_ln703_147_reg_1304 - data_12_V_read13_reg_1156_pp0_iter2_reg);

assign sub_ln703_24_fu_502_p2 = (add_ln703_150_fu_476_p2 - data_12_V_read13_reg_1156_pp0_iter2_reg);

assign sub_ln703_25_fu_517_p2 = (add_ln703_152_fu_493_p2 - data_13_V_read14_reg_1147_pp0_iter2_reg);

assign sub_ln703_26_fu_527_p2 = (add_ln703_153_fu_507_p2 - data_13_V_read14_reg_1147_pp0_iter2_reg);

assign sub_ln703_27_fu_532_p2 = (add_ln703_154_fu_512_p2 - data_13_V_read14_reg_1147_pp0_iter2_reg);

assign sub_ln703_28_fu_537_p2 = (add_ln703_155_fu_522_p2 - data_14_V_read15_reg_1138_pp0_iter2_reg);

assign sub_ln703_29_fu_575_p2 = (sub_ln703_26_reg_1324 - data_14_V_read15_reg_1138_pp0_iter3_reg);

assign sub_ln703_2_fu_292_p2 = (data_2_V_read_8_reg_1240 - add_ln703_reg_1246);

assign sub_ln703_30_fu_542_p2 = (sub_ln703_27_fu_532_p2 - data_14_V_read15_reg_1138_pp0_iter2_reg);

assign sub_ln703_31_fu_579_p2 = (add_ln703_156_fu_571_p2 - data_15_V_read16_reg_1129_pp0_iter3_reg);

assign sub_ln703_32_fu_584_p2 = (sub_ln703_28_reg_1329 - data_15_V_read16_reg_1129_pp0_iter3_reg);

assign sub_ln703_33_fu_562_p2 = (add_ln703_159_fu_556_p2 - data_16_V_read_7_reg_1120_pp0_iter2_reg);

assign sub_ln703_34_fu_597_p2 = (sub_ln703_32_fu_584_p2 - data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign sub_ln703_35_fu_602_p2 = (add_ln703_160_fu_588_p2 - data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign sub_ln703_36_fu_607_p2 = (add_ln703_161_fu_593_p2 - data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign sub_ln703_37_fu_612_p2 = (sub_ln703_33_reg_1339 - data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign sub_ln703_38_fu_626_p2 = (add_ln703_162_fu_616_p2 - data_18_V_read_6_reg_1103_pp0_iter3_reg);

assign sub_ln703_39_fu_666_p2 = (add_ln703_163_reg_1350 - data_18_V_read_6_reg_1103_pp0_iter4_reg);

assign sub_ln703_3_fu_296_p2 = (sub_ln703_1_reg_1252 - data_3_V_read_8_reg_1232);

assign sub_ln703_40_fu_670_p2 = (sub_ln703_38_reg_1355 - data_19_V_read_6_reg_1095_pp0_iter4_reg);

assign sub_ln703_41_fu_646_p2 = (add_ln703_165_fu_635_p2 - data_19_V_read_6_reg_1095_pp0_iter3_reg);

assign sub_ln703_42_fu_679_p2 = (add_ln703_167_reg_1360 - data_20_V_read21_reg_1086_pp0_iter4_reg);

assign sub_ln703_43_fu_683_p2 = (add_ln703_168_fu_674_p2 - data_20_V_read21_reg_1086_pp0_iter4_reg);

assign sub_ln703_44_fu_688_p2 = (sub_ln703_41_reg_1365 - data_20_V_read21_reg_1086_pp0_iter4_reg);

assign sub_ln703_45_fu_692_p2 = (sub_ln703_42_fu_679_p2 - data_21_V_read22_reg_1077_pp0_iter4_reg);

assign sub_ln703_46_fu_697_p2 = (sub_ln703_43_fu_683_p2 - data_21_V_read22_reg_1077_pp0_iter4_reg);

assign sub_ln703_47_fu_707_p2 = (sub_ln703_45_fu_692_p2 - data_22_V_read23_reg_1068_pp0_iter4_reg);

assign sub_ln703_48_fu_727_p2 = (add_ln703_169_fu_702_p2 - data_22_V_read23_reg_1068_pp0_iter4_reg);

assign sub_ln703_49_fu_737_p2 = (add_ln703_172_fu_721_p2 - data_23_V_read24_reg_1059_pp0_iter4_reg);

assign sub_ln703_4_fu_309_p2 = (sub_ln703_2_fu_292_p2 - data_3_V_read_8_reg_1232);

assign sub_ln703_50_fu_742_p2 = (sub_ln703_48_fu_727_p2 - data_23_V_read24_reg_1059_pp0_iter4_reg);

assign sub_ln703_51_fu_779_p2 = (add_ln703_173_reg_1380 - data_24_V_read25_reg_1050_pp0_iter5_reg);

assign sub_ln703_52_fu_783_p2 = (sub_ln703_49_reg_1385 - data_24_V_read25_reg_1050_pp0_iter5_reg);

assign sub_ln703_53_fu_787_p2 = (sub_ln703_50_reg_1390 - data_24_V_read25_reg_1050_pp0_iter5_reg);

assign sub_ln703_54_fu_791_p2 = (add_ln703_181_fu_775_p2 - data_25_V_read26_reg_1041_pp0_iter5_reg);

assign sub_ln703_55_fu_796_p2 = (sub_ln703_51_fu_779_p2 - data_25_V_read26_reg_1041_pp0_iter5_reg);

assign sub_ln703_56_fu_801_p2 = (sub_ln703_52_fu_783_p2 - data_25_V_read26_reg_1041_pp0_iter5_reg);

assign sub_ln703_57_fu_820_p2 = (sub_ln703_54_fu_791_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_58_fu_825_p2 = (sub_ln703_56_fu_801_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_59_fu_830_p2 = (add_ln703_185_fu_810_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_5_fu_319_p2 = (add_ln703_131_fu_304_p2 - data_4_V_read_8_reg_1224);

assign sub_ln703_60_fu_835_p2 = (add_ln703_186_fu_815_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_61_fu_840_p2 = (sub_ln703_57_fu_820_p2 - data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign sub_ln703_62_fu_860_p2 = (sub_ln703_60_fu_835_p2 - data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign sub_ln703_63_fu_879_p2 = (sub_ln703_61_reg_1405 - data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign sub_ln703_64_fu_865_p2 = (add_ln703_188_fu_849_p2 - data_28_V_read_6_reg_1014_pp0_iter5_reg);

assign sub_ln703_65_fu_883_p2 = (add_ln703_189_reg_1410 - data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign sub_ln703_66_fu_891_p2 = (sub_ln703_63_fu_879_p2 - data_29_V_read_6_reg_1006_pp0_iter6_reg);

assign sub_ln703_67_fu_901_p2 = (add_ln703_190_fu_887_p2 - data_29_V_read_6_reg_1006_pp0_iter6_reg);

assign sub_ln703_68_fu_906_p2 = (sub_ln703_66_fu_891_p2 - data_30_V_read31_reg_998_pp0_iter6_reg);

assign sub_ln703_69_fu_924_p2 = (add_ln703_191_fu_896_p2 - data_30_V_read31_reg_998_pp0_iter6_reg);

assign sub_ln703_6_fu_324_p2 = (sub_ln703_4_fu_309_p2 - data_4_V_read_8_reg_1224);

assign sub_ln703_70_fu_929_p2 = (sub_ln703_68_fu_906_p2 - data_31_V_read32_reg_989_pp0_iter6_reg);

assign sub_ln703_7_fu_373_p2 = (sub_ln703_5_reg_1258 - data_5_V_read_7_reg_1215_pp0_iter1_reg);

assign sub_ln703_8_fu_329_p2 = (add_ln703_132_fu_314_p2 - data_5_V_read_7_reg_1215);

assign sub_ln703_9_fu_353_p2 = (sub_ln703_8_fu_329_p2 - data_6_V_read_7_reg_1208);

assign sub_ln703_fu_274_p2 = (data_0_V_read_int_reg - data_1_V_read_int_reg);

endmodule //dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0
// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2019.2 (64-bit)
// Copyright 1986-2019 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module myproject_mul_16s_10ns_26_2_0_MulnS_4(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [10 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
`timescale 1 ns / 1 ps
module myproject_mul_16s_10ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_10ns_26_2_0_MulnS_4 myproject_mul_16s_10ns_26_2_0_MulnS_4_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2019.2 (64-bit)
// Copyright 1986-2019 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module myproject_mul_16s_11ns_26_2_0_MulnS_1(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [11 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
`timescale 1 ns / 1 ps
module myproject_mul_16s_11ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_11ns_26_2_0_MulnS_1 myproject_mul_16s_11ns_26_2_0_MulnS_1_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2019.2 (64-bit)
// Copyright 1986-2019 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module myproject_mul_16s_12ns_26_2_0_MulnS_0(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [12 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
`timescale 1 ns / 1 ps
module myproject_mul_16s_12ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_12ns_26_2_0_MulnS_0 myproject_mul_16s_12ns_26_2_0_MulnS_0_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2019.2 (64-bit)
// Copyright 1986-2019 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module myproject_mul_16s_13ns_26_2_0_MulnS_2(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [13 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
`timescale 1 ns / 1 ps
module myproject_mul_16s_13ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_13ns_26_2_0_MulnS_2 myproject_mul_16s_13ns_26_2_0_MulnS_2_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2019.2 (64-bit)
// Copyright 1986-2019 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module myproject_mul_16s_8ns_24_2_0_MulnS_5(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [8 - 1 : 0] b;
output[24 - 1 : 0] p;
reg  [24 - 1 : 0] p;
wire  [24 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
`timescale 1 ns / 1 ps
module myproject_mul_16s_8ns_24_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_8ns_24_2_0_MulnS_5 myproject_mul_16s_8ns_24_2_0_MulnS_5_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

// ==============================================================
// Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC v2019.2 (64-bit)
// Copyright 1986-2019 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module myproject_mul_16s_9ns_25_2_0_MulnS_3(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [9 - 1 : 0] b;
output[25 - 1 : 0] p;
reg  [25 - 1 : 0] p;
wire  [25 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
`timescale 1 ns / 1 ps
module myproject_mul_16s_9ns_25_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_9ns_25_2_0_MulnS_3 myproject_mul_16s_9ns_25_2_0_MulnS_3_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 


module myproject (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        input1_V_ap_vld,
        input1_V,
        layer16_out_0_V,
        layer16_out_0_V_ap_vld,
        layer16_out_1_V,
        layer16_out_1_V_ap_vld,
        layer16_out_2_V,
        layer16_out_2_V_ap_vld,
        layer16_out_3_V,
        layer16_out_3_V_ap_vld,
        layer16_out_4_V,
        layer16_out_4_V_ap_vld,
        const_size_in_1,
        const_size_in_1_ap_vld,
        const_size_out_1,
        const_size_out_1_ap_vld
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input   input1_V_ap_vld;
input  [255:0] input1_V;
output  [15:0] layer16_out_0_V;
output   layer16_out_0_V_ap_vld;
output  [15:0] layer16_out_1_V;
output   layer16_out_1_V_ap_vld;
output  [15:0] layer16_out_2_V;
output   layer16_out_2_V_ap_vld;
output  [15:0] layer16_out_3_V;
output   layer16_out_3_V_ap_vld;
output  [15:0] layer16_out_4_V;
output   layer16_out_4_V_ap_vld;
output  [15:0] const_size_in_1;
output   const_size_in_1_ap_vld;
output  [15:0] const_size_out_1;
output   const_size_out_1_ap_vld;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg layer16_out_0_V_ap_vld;
reg layer16_out_1_V_ap_vld;
reg layer16_out_2_V_ap_vld;
reg layer16_out_3_V_ap_vld;
reg layer16_out_4_V_ap_vld;
reg const_size_in_1_ap_vld;
reg const_size_out_1_ap_vld;

reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
reg    ap_enable_reg_pp0_iter23;
reg    ap_enable_reg_pp0_iter24;
reg    ap_enable_reg_pp0_iter25;
reg    ap_enable_reg_pp0_iter26;
reg    ap_enable_reg_pp0_iter27;
reg    ap_enable_reg_pp0_iter28;
reg    ap_enable_reg_pp0_iter29;
reg    ap_enable_reg_pp0_iter30;
reg    ap_enable_reg_pp0_iter31;
reg    ap_enable_reg_pp0_iter32;
reg    ap_enable_reg_pp0_iter33;
reg    ap_enable_reg_pp0_iter34;
reg    ap_enable_reg_pp0_iter35;
reg    ap_enable_reg_pp0_iter36;
reg    ap_enable_reg_pp0_iter37;
reg    ap_enable_reg_pp0_iter38;
reg    ap_enable_reg_pp0_iter39;
reg    ap_enable_reg_pp0_iter40;
reg    ap_enable_reg_pp0_iter41;
reg    ap_enable_reg_pp0_iter42;
reg    ap_enable_reg_pp0_iter43;
reg    ap_enable_reg_pp0_iter44;
reg    ap_enable_reg_pp0_iter45;
reg    ap_enable_reg_pp0_iter46;
reg    ap_enable_reg_pp0_iter47;
reg    ap_enable_reg_pp0_iter48;
reg    ap_enable_reg_pp0_iter49;
reg    ap_enable_reg_pp0_iter50;
reg    ap_enable_reg_pp0_iter51;
reg    ap_enable_reg_pp0_iter52;
reg    ap_enable_reg_pp0_iter53;
reg    ap_enable_reg_pp0_iter54;
reg    ap_enable_reg_pp0_iter55;
reg    ap_enable_reg_pp0_iter56;
reg    ap_enable_reg_pp0_iter57;
reg    ap_enable_reg_pp0_iter58;
reg    ap_enable_reg_pp0_iter59;
reg    ap_enable_reg_pp0_iter60;
reg    ap_enable_reg_pp0_iter61;
reg    ap_enable_reg_pp0_iter62;
reg    ap_enable_reg_pp0_iter63;
reg    ap_enable_reg_pp0_iter64;
reg    ap_enable_reg_pp0_iter65;
reg    ap_enable_reg_pp0_iter66;
reg    ap_enable_reg_pp0_iter67;
reg    ap_idle_pp0;
reg    input1_V_ap_vld_in_sig;
reg    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_state19_pp0_stage0_iter18;
wire    ap_block_state20_pp0_stage0_iter19;
wire    ap_block_state21_pp0_stage0_iter20;
wire    ap_block_state22_pp0_stage0_iter21;
wire    ap_block_state23_pp0_stage0_iter22;
wire    ap_block_state24_pp0_stage0_iter23;
wire    ap_block_state25_pp0_stage0_iter24;
wire    ap_block_state26_pp0_stage0_iter25;
wire    ap_block_state27_pp0_stage0_iter26;
wire    ap_block_state28_pp0_stage0_iter27;
wire    ap_block_state29_pp0_stage0_iter28;
wire    ap_block_state30_pp0_stage0_iter29;
wire    ap_block_state31_pp0_stage0_iter30;
wire    ap_block_state32_pp0_stage0_iter31;
wire    ap_block_state33_pp0_stage0_iter32;
wire    ap_block_state34_pp0_stage0_iter33;
wire    ap_block_state35_pp0_stage0_iter34;
wire    ap_block_state36_pp0_stage0_iter35;
wire    ap_block_state37_pp0_stage0_iter36;
wire    ap_block_state38_pp0_stage0_iter37;
wire    ap_block_state39_pp0_stage0_iter38;
wire    ap_block_state40_pp0_stage0_iter39;
wire    ap_block_state41_pp0_stage0_iter40;
wire    ap_block_state42_pp0_stage0_iter41;
wire    ap_block_state43_pp0_stage0_iter42;
wire    ap_block_state44_pp0_stage0_iter43;
wire    ap_block_state45_pp0_stage0_iter44;
wire    ap_block_state46_pp0_stage0_iter45;
wire    ap_block_state47_pp0_stage0_iter46;
wire    ap_block_state48_pp0_stage0_iter47;
wire    ap_block_state49_pp0_stage0_iter48;
wire    ap_block_state50_pp0_stage0_iter49;
wire    ap_block_state51_pp0_stage0_iter50;
wire    ap_block_state52_pp0_stage0_iter51;
wire    ap_block_state53_pp0_stage0_iter52;
wire    ap_block_state54_pp0_stage0_iter53;
wire    ap_block_state55_pp0_stage0_iter54;
wire    ap_block_state56_pp0_stage0_iter55;
wire    ap_block_state57_pp0_stage0_iter56;
wire    ap_block_state58_pp0_stage0_iter57;
wire    ap_block_state59_pp0_stage0_iter58;
wire    ap_block_state60_pp0_stage0_iter59;
wire    ap_block_state61_pp0_stage0_iter60;
wire    ap_block_state62_pp0_stage0_iter61;
wire    ap_block_state63_pp0_stage0_iter62;
wire    ap_block_state64_pp0_stage0_iter63;
wire    ap_block_state65_pp0_stage0_iter64;
wire    ap_block_state66_pp0_stage0_iter65;
wire    ap_block_state67_pp0_stage0_iter66;
wire    ap_block_state68_pp0_stage0_iter67;
reg    ap_block_pp0_stage0_11001;
reg   [255:0] input1_V_preg;
reg   [255:0] input1_V_in_sig;
reg    input1_V_ap_vld_preg;
reg    input1_V_blk_n;
wire    ap_block_pp0_stage0;
reg   [15:0] layer2_out_0_V_reg_2146;
reg   [15:0] layer2_out_1_V_reg_2151;
reg   [15:0] layer2_out_2_V_reg_2156;
reg   [15:0] layer2_out_3_V_reg_2161;
reg   [15:0] layer2_out_4_V_reg_2166;
reg   [15:0] layer2_out_5_V_reg_2171;
reg   [15:0] layer2_out_6_V_reg_2176;
reg   [15:0] layer2_out_7_V_reg_2181;
reg   [15:0] layer2_out_8_V_reg_2186;
reg   [15:0] layer2_out_9_V_reg_2191;
reg   [15:0] layer2_out_10_V_reg_2196;
reg   [15:0] layer2_out_11_V_reg_2201;
reg   [15:0] layer2_out_12_V_reg_2206;
reg   [15:0] layer2_out_13_V_reg_2211;
reg   [15:0] layer2_out_14_V_reg_2216;
reg   [15:0] layer2_out_15_V_reg_2221;
reg   [15:0] layer2_out_16_V_reg_2226;
reg   [15:0] layer2_out_17_V_reg_2231;
reg   [15:0] layer2_out_18_V_reg_2236;
reg   [15:0] layer2_out_19_V_reg_2241;
reg   [15:0] layer2_out_20_V_reg_2246;
reg   [15:0] layer2_out_21_V_reg_2251;
reg   [15:0] layer2_out_22_V_reg_2256;
reg   [15:0] layer2_out_23_V_reg_2261;
reg   [15:0] layer2_out_24_V_reg_2266;
reg   [15:0] layer2_out_25_V_reg_2271;
reg   [15:0] layer2_out_26_V_reg_2276;
reg   [15:0] layer2_out_27_V_reg_2281;
reg   [15:0] layer2_out_28_V_reg_2286;
reg   [15:0] layer2_out_29_V_reg_2291;
reg   [15:0] layer2_out_30_V_reg_2296;
reg   [15:0] layer2_out_31_V_reg_2301;
reg   [15:0] layer2_out_32_V_reg_2306;
reg   [15:0] layer2_out_33_V_reg_2311;
reg   [15:0] layer2_out_34_V_reg_2316;
reg   [15:0] layer2_out_35_V_reg_2321;
reg   [15:0] layer2_out_36_V_reg_2326;
reg   [15:0] layer2_out_37_V_reg_2331;
reg   [15:0] layer2_out_38_V_reg_2336;
reg   [15:0] layer2_out_39_V_reg_2341;
reg   [15:0] layer2_out_40_V_reg_2346;
reg   [15:0] layer2_out_41_V_reg_2351;
reg   [15:0] layer2_out_42_V_reg_2356;
reg   [15:0] layer2_out_43_V_reg_2361;
reg   [15:0] layer2_out_44_V_reg_2366;
reg   [15:0] layer2_out_45_V_reg_2371;
reg   [15:0] layer2_out_46_V_reg_2376;
reg   [15:0] layer2_out_47_V_reg_2381;
reg   [15:0] layer2_out_48_V_reg_2386;
reg   [15:0] layer2_out_49_V_reg_2391;
reg   [15:0] layer2_out_50_V_reg_2396;
reg   [15:0] layer2_out_51_V_reg_2401;
reg   [15:0] layer2_out_52_V_reg_2406;
reg   [15:0] layer2_out_53_V_reg_2411;
reg   [15:0] layer2_out_54_V_reg_2416;
reg   [15:0] layer2_out_55_V_reg_2421;
reg   [15:0] layer2_out_56_V_reg_2426;
reg   [15:0] layer2_out_57_V_reg_2431;
reg   [15:0] layer2_out_58_V_reg_2436;
reg   [15:0] layer2_out_59_V_reg_2441;
reg   [15:0] layer2_out_60_V_reg_2446;
reg   [15:0] layer2_out_61_V_reg_2451;
reg   [15:0] layer2_out_62_V_reg_2456;
reg   [15:0] layer2_out_63_V_reg_2461;
reg   [15:0] layer4_out_0_V_reg_2466;
reg   [15:0] layer4_out_1_V_reg_2471;
reg   [15:0] layer4_out_2_V_reg_2476;
reg   [15:0] layer4_out_3_V_reg_2481;
reg   [15:0] layer4_out_4_V_reg_2486;
reg   [15:0] layer4_out_5_V_reg_2491;
reg   [15:0] layer4_out_6_V_reg_2496;
reg   [15:0] layer4_out_7_V_reg_2501;
reg   [15:0] layer4_out_8_V_reg_2506;
reg   [15:0] layer4_out_9_V_reg_2511;
reg   [15:0] layer4_out_10_V_reg_2516;
reg   [15:0] layer4_out_11_V_reg_2521;
reg   [15:0] layer4_out_12_V_reg_2526;
reg   [15:0] layer4_out_13_V_reg_2531;
reg   [15:0] layer4_out_14_V_reg_2536;
reg   [15:0] layer4_out_15_V_reg_2541;
reg   [15:0] layer4_out_16_V_reg_2546;
reg   [15:0] layer4_out_17_V_reg_2551;
reg   [15:0] layer4_out_18_V_reg_2556;
reg   [15:0] layer4_out_19_V_reg_2561;
reg   [15:0] layer4_out_20_V_reg_2566;
reg   [15:0] layer4_out_21_V_reg_2571;
reg   [15:0] layer4_out_22_V_reg_2576;
reg   [15:0] layer4_out_23_V_reg_2581;
reg   [15:0] layer4_out_24_V_reg_2586;
reg   [15:0] layer4_out_25_V_reg_2591;
reg   [15:0] layer4_out_26_V_reg_2596;
reg   [15:0] layer4_out_27_V_reg_2601;
reg   [15:0] layer4_out_28_V_reg_2606;
reg   [15:0] layer4_out_29_V_reg_2611;
reg   [15:0] layer4_out_30_V_reg_2616;
reg   [15:0] layer4_out_31_V_reg_2621;
reg   [15:0] layer4_out_32_V_reg_2626;
reg   [15:0] layer4_out_33_V_reg_2631;
reg   [15:0] layer4_out_34_V_reg_2636;
reg   [15:0] layer4_out_35_V_reg_2641;
reg   [15:0] layer4_out_36_V_reg_2646;
reg   [15:0] layer4_out_37_V_reg_2651;
reg   [15:0] layer4_out_38_V_reg_2656;
reg   [15:0] layer4_out_39_V_reg_2661;
reg   [15:0] layer4_out_40_V_reg_2666;
reg   [15:0] layer4_out_41_V_reg_2671;
reg   [15:0] layer4_out_42_V_reg_2676;
reg   [15:0] layer4_out_43_V_reg_2681;
reg   [15:0] layer4_out_44_V_reg_2686;
reg   [15:0] layer4_out_45_V_reg_2691;
reg   [15:0] layer4_out_46_V_reg_2696;
reg   [15:0] layer4_out_47_V_reg_2701;
reg   [15:0] layer4_out_48_V_reg_2706;
reg   [15:0] layer4_out_49_V_reg_2711;
reg   [15:0] layer4_out_50_V_reg_2716;
reg   [15:0] layer4_out_51_V_reg_2721;
reg   [15:0] layer4_out_52_V_reg_2726;
reg   [15:0] layer4_out_53_V_reg_2731;
reg   [15:0] layer4_out_54_V_reg_2736;
reg   [15:0] layer4_out_55_V_reg_2741;
reg   [15:0] layer4_out_56_V_reg_2746;
reg   [15:0] layer4_out_57_V_reg_2751;
reg   [15:0] layer4_out_58_V_reg_2756;
reg   [15:0] layer4_out_59_V_reg_2761;
reg   [15:0] layer4_out_60_V_reg_2766;
reg   [15:0] layer4_out_61_V_reg_2771;
reg   [15:0] layer4_out_62_V_reg_2776;
reg   [15:0] layer4_out_63_V_reg_2781;
reg   [15:0] layer5_out_0_V_reg_2786;
reg   [15:0] layer5_out_1_V_reg_2791;
reg   [15:0] layer5_out_2_V_reg_2796;
reg   [15:0] layer5_out_3_V_reg_2801;
reg   [15:0] layer5_out_4_V_reg_2806;
reg   [15:0] layer5_out_5_V_reg_2811;
reg   [15:0] layer5_out_6_V_reg_2816;
reg   [15:0] layer5_out_7_V_reg_2821;
reg   [15:0] layer5_out_8_V_reg_2826;
reg   [15:0] layer5_out_9_V_reg_2831;
reg   [15:0] layer5_out_10_V_reg_2836;
reg   [15:0] layer5_out_11_V_reg_2841;
reg   [15:0] layer5_out_12_V_reg_2846;
reg   [15:0] layer5_out_13_V_reg_2851;
reg   [15:0] layer5_out_14_V_reg_2856;
reg   [15:0] layer5_out_15_V_reg_2861;
reg   [15:0] layer5_out_16_V_reg_2866;
reg   [15:0] layer5_out_17_V_reg_2871;
reg   [15:0] layer5_out_18_V_reg_2876;
reg   [15:0] layer5_out_19_V_reg_2881;
reg   [15:0] layer5_out_20_V_reg_2886;
reg   [15:0] layer5_out_21_V_reg_2891;
reg   [15:0] layer5_out_22_V_reg_2896;
reg   [15:0] layer5_out_23_V_reg_2901;
reg   [15:0] layer5_out_24_V_reg_2906;
reg   [15:0] layer5_out_25_V_reg_2911;
reg   [15:0] layer5_out_26_V_reg_2916;
reg   [15:0] layer5_out_27_V_reg_2921;
reg   [15:0] layer5_out_28_V_reg_2926;
reg   [15:0] layer5_out_29_V_reg_2931;
reg   [15:0] layer5_out_30_V_reg_2936;
reg   [15:0] layer5_out_31_V_reg_2941;
reg   [15:0] layer5_out_32_V_reg_2946;
reg   [15:0] layer5_out_33_V_reg_2951;
reg   [15:0] layer5_out_34_V_reg_2956;
reg   [15:0] layer5_out_35_V_reg_2961;
reg   [15:0] layer5_out_36_V_reg_2966;
reg   [15:0] layer5_out_37_V_reg_2971;
reg   [15:0] layer5_out_38_V_reg_2976;
reg   [15:0] layer5_out_39_V_reg_2981;
reg   [15:0] layer5_out_40_V_reg_2986;
reg   [15:0] layer5_out_41_V_reg_2991;
reg   [15:0] layer5_out_42_V_reg_2996;
reg   [15:0] layer5_out_43_V_reg_3001;
reg   [15:0] layer5_out_44_V_reg_3006;
reg   [15:0] layer5_out_45_V_reg_3011;
reg   [15:0] layer5_out_46_V_reg_3016;
reg   [15:0] layer5_out_47_V_reg_3021;
reg   [15:0] layer5_out_48_V_reg_3026;
reg   [15:0] layer5_out_49_V_reg_3031;
reg   [15:0] layer5_out_50_V_reg_3036;
reg   [15:0] layer5_out_51_V_reg_3041;
reg   [15:0] layer5_out_52_V_reg_3046;
reg   [15:0] layer5_out_53_V_reg_3051;
reg   [15:0] layer5_out_54_V_reg_3056;
reg   [15:0] layer5_out_55_V_reg_3061;
reg   [15:0] layer5_out_56_V_reg_3066;
reg   [15:0] layer5_out_57_V_reg_3071;
reg   [15:0] layer5_out_58_V_reg_3076;
reg   [15:0] layer5_out_59_V_reg_3081;
reg   [15:0] layer5_out_60_V_reg_3086;
reg   [15:0] layer5_out_61_V_reg_3091;
reg   [15:0] layer5_out_62_V_reg_3096;
reg   [15:0] layer5_out_63_V_reg_3101;
reg   [15:0] layer6_out_0_V_reg_3106;
reg   [15:0] layer6_out_1_V_reg_3111;
reg   [15:0] layer6_out_2_V_reg_3116;
reg   [15:0] layer6_out_3_V_reg_3121;
reg   [15:0] layer6_out_4_V_reg_3126;
reg   [15:0] layer6_out_5_V_reg_3131;
reg   [15:0] layer6_out_6_V_reg_3136;
reg   [15:0] layer6_out_7_V_reg_3141;
reg   [15:0] layer6_out_8_V_reg_3146;
reg   [15:0] layer6_out_9_V_reg_3151;
reg   [15:0] layer6_out_10_V_reg_3156;
reg   [15:0] layer6_out_11_V_reg_3161;
reg   [15:0] layer6_out_12_V_reg_3166;
reg   [15:0] layer6_out_13_V_reg_3171;
reg   [15:0] layer6_out_14_V_reg_3176;
reg   [15:0] layer6_out_15_V_reg_3181;
reg   [15:0] layer6_out_16_V_reg_3186;
reg   [15:0] layer6_out_17_V_reg_3191;
reg   [15:0] layer6_out_18_V_reg_3196;
reg   [15:0] layer6_out_19_V_reg_3201;
reg   [15:0] layer6_out_20_V_reg_3206;
reg   [15:0] layer6_out_21_V_reg_3211;
reg   [15:0] layer6_out_22_V_reg_3216;
reg   [15:0] layer6_out_23_V_reg_3221;
reg   [15:0] layer6_out_24_V_reg_3226;
reg   [15:0] layer6_out_25_V_reg_3231;
reg   [15:0] layer6_out_26_V_reg_3236;
reg   [15:0] layer6_out_27_V_reg_3241;
reg   [15:0] layer6_out_28_V_reg_3246;
reg   [15:0] layer6_out_29_V_reg_3251;
reg   [15:0] layer6_out_30_V_reg_3256;
reg   [15:0] layer6_out_31_V_reg_3261;
reg   [15:0] layer8_out_0_V_reg_3266;
reg   [15:0] layer8_out_1_V_reg_3271;
reg   [15:0] layer8_out_2_V_reg_3276;
reg   [15:0] layer8_out_3_V_reg_3281;
reg   [15:0] layer8_out_4_V_reg_3286;
reg   [15:0] layer8_out_5_V_reg_3291;
reg   [15:0] layer8_out_6_V_reg_3296;
reg   [15:0] layer8_out_7_V_reg_3301;
reg   [15:0] layer8_out_8_V_reg_3306;
reg   [15:0] layer8_out_9_V_reg_3311;
reg   [15:0] layer8_out_10_V_reg_3316;
reg   [15:0] layer8_out_11_V_reg_3321;
reg   [15:0] layer8_out_12_V_reg_3326;
reg   [15:0] layer8_out_13_V_reg_3331;
reg   [15:0] layer8_out_14_V_reg_3336;
reg   [15:0] layer8_out_15_V_reg_3341;
reg   [15:0] layer8_out_16_V_reg_3346;
reg   [15:0] layer8_out_17_V_reg_3351;
reg   [15:0] layer8_out_18_V_reg_3356;
reg   [15:0] layer8_out_19_V_reg_3361;
reg   [15:0] layer8_out_20_V_reg_3366;
reg   [15:0] layer8_out_21_V_reg_3371;
reg   [15:0] layer8_out_22_V_reg_3376;
reg   [15:0] layer8_out_23_V_reg_3381;
reg   [15:0] layer8_out_24_V_reg_3386;
reg   [15:0] layer8_out_25_V_reg_3391;
reg   [15:0] layer8_out_26_V_reg_3396;
reg   [15:0] layer8_out_27_V_reg_3401;
reg   [15:0] layer8_out_28_V_reg_3406;
reg   [15:0] layer8_out_29_V_reg_3411;
reg   [15:0] layer8_out_30_V_reg_3416;
reg   [15:0] layer8_out_31_V_reg_3421;
reg   [15:0] layer9_out_0_V_reg_3426;
reg   [15:0] layer9_out_1_V_reg_3431;
reg   [15:0] layer9_out_2_V_reg_3436;
reg   [15:0] layer9_out_3_V_reg_3441;
reg   [15:0] layer9_out_4_V_reg_3446;
reg   [15:0] layer9_out_5_V_reg_3451;
reg   [15:0] layer9_out_6_V_reg_3456;
reg   [15:0] layer9_out_7_V_reg_3461;
reg   [15:0] layer9_out_8_V_reg_3466;
reg   [15:0] layer9_out_9_V_reg_3471;
reg   [15:0] layer9_out_10_V_reg_3476;
reg   [15:0] layer9_out_11_V_reg_3481;
reg   [15:0] layer9_out_12_V_reg_3486;
reg   [15:0] layer9_out_13_V_reg_3491;
reg   [15:0] layer9_out_14_V_reg_3496;
reg   [15:0] layer9_out_15_V_reg_3501;
reg   [15:0] layer9_out_16_V_reg_3506;
reg   [15:0] layer9_out_17_V_reg_3511;
reg   [15:0] layer9_out_18_V_reg_3516;
reg   [15:0] layer9_out_19_V_reg_3521;
reg   [15:0] layer9_out_20_V_reg_3526;
reg   [15:0] layer9_out_21_V_reg_3531;
reg   [15:0] layer9_out_22_V_reg_3536;
reg   [15:0] layer9_out_23_V_reg_3541;
reg   [15:0] layer9_out_24_V_reg_3546;
reg   [15:0] layer9_out_25_V_reg_3551;
reg   [15:0] layer9_out_26_V_reg_3556;
reg   [15:0] layer9_out_27_V_reg_3561;
reg   [15:0] layer9_out_28_V_reg_3566;
reg   [15:0] layer9_out_29_V_reg_3571;
reg   [15:0] layer9_out_30_V_reg_3576;
reg   [15:0] layer9_out_31_V_reg_3581;
reg   [15:0] layer10_out_0_V_reg_3586;
reg   [15:0] layer10_out_1_V_reg_3591;
reg   [15:0] layer10_out_2_V_reg_3596;
reg   [15:0] layer10_out_3_V_reg_3601;
reg   [15:0] layer10_out_4_V_reg_3606;
reg   [15:0] layer10_out_5_V_reg_3611;
reg   [15:0] layer10_out_6_V_reg_3616;
reg   [15:0] layer10_out_7_V_reg_3621;
reg   [15:0] layer10_out_8_V_reg_3626;
reg   [15:0] layer10_out_9_V_reg_3631;
reg   [15:0] layer10_out_10_V_reg_3636;
reg   [15:0] layer10_out_11_V_reg_3641;
reg   [15:0] layer10_out_12_V_reg_3646;
reg   [15:0] layer10_out_13_V_reg_3651;
reg   [15:0] layer10_out_14_V_reg_3656;
reg   [15:0] layer10_out_15_V_reg_3661;
reg   [15:0] layer10_out_16_V_reg_3666;
reg   [15:0] layer10_out_17_V_reg_3671;
reg   [15:0] layer10_out_18_V_reg_3676;
reg   [15:0] layer10_out_19_V_reg_3681;
reg   [15:0] layer10_out_20_V_reg_3686;
reg   [15:0] layer10_out_21_V_reg_3691;
reg   [15:0] layer10_out_22_V_reg_3696;
reg   [15:0] layer10_out_23_V_reg_3701;
reg   [15:0] layer10_out_24_V_reg_3706;
reg   [15:0] layer10_out_25_V_reg_3711;
reg   [15:0] layer10_out_26_V_reg_3716;
reg   [15:0] layer10_out_27_V_reg_3721;
reg   [15:0] layer10_out_28_V_reg_3726;
reg   [15:0] layer10_out_29_V_reg_3731;
reg   [15:0] layer10_out_30_V_reg_3736;
reg   [15:0] layer10_out_31_V_reg_3741;
reg   [15:0] layer12_out_0_V_reg_3746;
reg   [15:0] layer12_out_1_V_reg_3751;
reg   [15:0] layer12_out_2_V_reg_3756;
reg   [15:0] layer12_out_3_V_reg_3761;
reg   [15:0] layer12_out_4_V_reg_3766;
reg   [15:0] layer12_out_5_V_reg_3771;
reg   [15:0] layer12_out_6_V_reg_3776;
reg   [15:0] layer12_out_7_V_reg_3781;
reg   [15:0] layer12_out_8_V_reg_3786;
reg   [15:0] layer12_out_9_V_reg_3791;
reg   [15:0] layer12_out_10_V_reg_3796;
reg   [15:0] layer12_out_11_V_reg_3801;
reg   [15:0] layer12_out_12_V_reg_3806;
reg   [15:0] layer12_out_13_V_reg_3811;
reg   [15:0] layer12_out_14_V_reg_3816;
reg   [15:0] layer12_out_15_V_reg_3821;
reg   [15:0] layer12_out_16_V_reg_3826;
reg   [15:0] layer12_out_17_V_reg_3831;
reg   [15:0] layer12_out_18_V_reg_3836;
reg   [15:0] layer12_out_19_V_reg_3841;
reg   [15:0] layer12_out_20_V_reg_3846;
reg   [15:0] layer12_out_21_V_reg_3851;
reg   [15:0] layer12_out_22_V_reg_3856;
reg   [15:0] layer12_out_23_V_reg_3861;
reg   [15:0] layer12_out_24_V_reg_3866;
reg   [15:0] layer12_out_25_V_reg_3871;
reg   [15:0] layer12_out_26_V_reg_3876;
reg   [15:0] layer12_out_27_V_reg_3881;
reg   [15:0] layer12_out_28_V_reg_3886;
reg   [15:0] layer12_out_29_V_reg_3891;
reg   [15:0] layer12_out_30_V_reg_3896;
reg   [15:0] layer12_out_31_V_reg_3901;
reg   [15:0] layer13_out_0_V_reg_3906;
reg   [15:0] layer13_out_1_V_reg_3911;
reg   [15:0] layer13_out_2_V_reg_3916;
reg   [15:0] layer13_out_3_V_reg_3921;
reg   [15:0] layer13_out_4_V_reg_3926;
reg   [15:0] layer13_out_5_V_reg_3931;
reg   [15:0] layer13_out_6_V_reg_3936;
reg   [15:0] layer13_out_7_V_reg_3941;
reg   [15:0] layer13_out_8_V_reg_3946;
reg   [15:0] layer13_out_9_V_reg_3951;
reg   [15:0] layer13_out_10_V_reg_3956;
reg   [15:0] layer13_out_11_V_reg_3961;
reg   [15:0] layer13_out_12_V_reg_3966;
reg   [15:0] layer13_out_13_V_reg_3971;
reg   [15:0] layer13_out_14_V_reg_3976;
reg   [15:0] layer13_out_15_V_reg_3981;
reg   [15:0] layer13_out_16_V_reg_3986;
reg   [15:0] layer13_out_17_V_reg_3991;
reg   [15:0] layer13_out_18_V_reg_3996;
reg   [15:0] layer13_out_19_V_reg_4001;
reg   [15:0] layer13_out_20_V_reg_4006;
reg   [15:0] layer13_out_21_V_reg_4011;
reg   [15:0] layer13_out_22_V_reg_4016;
reg   [15:0] layer13_out_23_V_reg_4021;
reg   [15:0] layer13_out_24_V_reg_4026;
reg   [15:0] layer13_out_25_V_reg_4031;
reg   [15:0] layer13_out_26_V_reg_4036;
reg   [15:0] layer13_out_27_V_reg_4041;
reg   [15:0] layer13_out_28_V_reg_4046;
reg   [15:0] layer13_out_29_V_reg_4051;
reg   [15:0] layer13_out_30_V_reg_4056;
reg   [15:0] layer13_out_31_V_reg_4061;
reg   [15:0] layer14_out_0_V_reg_4066;
reg   [15:0] layer14_out_1_V_reg_4071;
reg   [15:0] layer14_out_2_V_reg_4076;
reg   [15:0] layer14_out_3_V_reg_4081;
reg   [15:0] layer14_out_4_V_reg_4086;
reg    ap_block_pp0_stage0_subdone;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_0;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_1;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_2;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_3;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_4;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_5;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_6;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_7;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_8;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_9;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_10;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_11;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_12;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_13;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_14;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_15;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_16;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_17;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_18;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_19;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_20;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_21;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_22;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_23;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_24;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_25;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_26;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_27;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_28;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_29;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_30;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_31;
reg    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call210;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call210;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call210;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call210;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call210;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call210;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call210;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call210;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call210;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call210;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call210;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call210;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call210;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call210;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call210;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call210;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call210;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call210;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call210;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call210;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call210;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call210;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call210;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call210;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call210;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call210;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call210;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call210;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call210;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call210;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call210;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call210;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call210;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call210;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call210;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call210;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call210;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call210;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call210;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call210;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call210;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call210;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call210;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call210;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call210;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call210;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call210;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call210;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call210;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call210;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call210;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call210;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call210;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call210;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call210;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call210;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call210;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call210;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call210;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call210;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call210;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call210;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call210;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call210;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call210;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call210;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call210;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call210;
reg    ap_block_pp0_stage0_11001_ignoreCallOp277;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_0;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_1;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_2;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_3;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_4;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_5;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_6;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_7;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_8;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_9;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_10;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_11;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_12;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_13;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_14;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_15;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_16;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_17;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_18;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_19;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_20;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_21;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_22;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_23;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_24;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_25;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_26;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_27;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_28;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_29;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_30;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_31;
reg    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call309;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call309;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call309;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call309;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call309;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call309;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call309;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call309;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call309;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call309;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call309;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call309;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call309;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call309;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call309;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call309;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call309;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call309;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call309;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call309;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call309;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call309;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call309;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call309;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call309;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call309;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call309;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call309;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call309;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call309;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call309;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call309;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call309;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call309;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call309;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call309;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call309;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call309;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call309;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call309;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call309;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call309;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call309;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call309;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call309;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call309;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call309;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call309;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call309;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call309;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call309;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call309;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call309;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call309;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call309;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call309;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call309;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call309;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call309;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call309;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call309;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call309;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call309;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call309;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call309;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call309;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call309;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call309;
reg    ap_block_pp0_stage0_11001_ignoreCallOp397;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_0;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_1;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_2;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_3;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_4;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_5;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_6;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_7;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_8;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_9;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_10;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_11;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_12;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_13;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_14;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_15;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_16;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_17;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_18;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_19;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_20;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_21;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_22;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_23;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_24;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_25;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_26;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_27;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_28;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_29;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_30;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_31;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_32;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_33;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_34;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_35;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_36;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_37;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_38;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_39;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_40;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_41;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_42;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_43;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_44;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_45;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_46;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_47;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_48;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_49;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_50;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_51;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_52;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_53;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_54;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_55;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_56;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_57;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_58;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_59;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_60;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_61;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_62;
wire   [15:0] grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_63;
reg    grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call15;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call15;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call15;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call15;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call15;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call15;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call15;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call15;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call15;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call15;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call15;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call15;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call15;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call15;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call15;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call15;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call15;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call15;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call15;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call15;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call15;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call15;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call15;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call15;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call15;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call15;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call15;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call15;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call15;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call15;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call15;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call15;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call15;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call15;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call15;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call15;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call15;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call15;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call15;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call15;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call15;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call15;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call15;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call15;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call15;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call15;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call15;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call15;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call15;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call15;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call15;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call15;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call15;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call15;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call15;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call15;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call15;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call15;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call15;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call15;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call15;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call15;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call15;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call15;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call15;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call15;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call15;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call15;
reg    ap_block_pp0_stage0_11001_ignoreCallOp70;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_0;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_1;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_2;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_3;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_4;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_5;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_6;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_7;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_8;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_9;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_10;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_11;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_12;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_13;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_14;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_15;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_16;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_17;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_18;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_19;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_20;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_21;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_22;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_23;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_24;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_25;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_26;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_27;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_28;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_29;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_30;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_31;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_32;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_33;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_34;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_35;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_36;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_37;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_38;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_39;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_40;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_41;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_42;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_43;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_44;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_45;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_46;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_47;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_48;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_49;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_50;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_51;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_52;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_53;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_54;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_55;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_56;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_57;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_58;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_59;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_60;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_61;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_62;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_63;
reg    grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call80;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call80;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call80;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call80;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call80;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call80;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call80;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call80;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call80;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call80;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call80;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call80;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call80;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call80;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call80;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call80;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call80;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call80;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call80;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call80;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call80;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call80;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call80;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call80;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call80;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call80;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call80;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call80;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call80;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call80;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call80;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call80;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call80;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call80;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call80;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call80;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call80;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call80;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call80;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call80;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call80;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call80;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call80;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call80;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call80;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call80;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call80;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call80;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call80;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call80;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call80;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call80;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call80;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call80;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call80;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call80;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call80;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call80;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call80;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call80;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call80;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call80;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call80;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call80;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call80;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call80;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call80;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call80;
reg    ap_block_pp0_stage0_11001_ignoreCallOp144;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_0;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_1;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_2;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_3;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_4;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_5;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_6;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_7;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_8;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_9;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_10;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_11;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_12;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_13;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_14;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_15;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_16;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_17;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_18;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_19;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_20;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_21;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_22;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_23;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_24;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_25;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_26;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_27;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_28;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_29;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_30;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_31;
reg    grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call342;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call342;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call342;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call342;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call342;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call342;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call342;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call342;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call342;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call342;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call342;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call342;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call342;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call342;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call342;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call342;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call342;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call342;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call342;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call342;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call342;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call342;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call342;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call342;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call342;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call342;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call342;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call342;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call342;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call342;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call342;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call342;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call342;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call342;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call342;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call342;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call342;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call342;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call342;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call342;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call342;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call342;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call342;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call342;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call342;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call342;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call342;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call342;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call342;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call342;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call342;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call342;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call342;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call342;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call342;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call342;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call342;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call342;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call342;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call342;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call342;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call342;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call342;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call342;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call342;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call342;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call342;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call342;
reg    ap_block_pp0_stage0_11001_ignoreCallOp440;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_0;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_1;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_2;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_3;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_4;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_5;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_6;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_7;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_8;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_9;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_10;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_11;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_12;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_13;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_14;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_15;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_16;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_17;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_18;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_19;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_20;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_21;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_22;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_23;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_24;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_25;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_26;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_27;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_28;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_29;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_30;
wire   [15:0] grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_31;
reg    grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call243;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call243;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call243;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call243;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call243;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call243;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call243;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call243;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call243;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call243;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call243;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call243;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call243;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call243;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call243;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call243;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call243;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call243;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call243;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call243;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call243;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call243;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call243;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call243;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call243;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call243;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call243;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call243;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call243;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call243;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call243;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call243;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call243;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call243;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call243;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call243;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call243;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call243;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call243;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call243;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call243;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call243;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call243;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call243;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call243;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call243;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call243;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call243;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call243;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call243;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call243;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call243;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call243;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call243;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call243;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call243;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call243;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call243;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call243;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call243;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call243;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call243;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call243;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call243;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call243;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call243;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call243;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call243;
reg    ap_block_pp0_stage0_11001_ignoreCallOp328;
wire   [15:0] grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_0;
wire   [15:0] grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_1;
wire   [15:0] grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_2;
wire   [15:0] grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_3;
wire   [15:0] grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_4;
reg    grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call408;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call408;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call408;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call408;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call408;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call408;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call408;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call408;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call408;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call408;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call408;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call408;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call408;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call408;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call408;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call408;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call408;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call408;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call408;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call408;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call408;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call408;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call408;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call408;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call408;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call408;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call408;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call408;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call408;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call408;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call408;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call408;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call408;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call408;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call408;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call408;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call408;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call408;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call408;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call408;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call408;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call408;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call408;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call408;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call408;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call408;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call408;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call408;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call408;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call408;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call408;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call408;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call408;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call408;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call408;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call408;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call408;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call408;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call408;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call408;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call408;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call408;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call408;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call408;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call408;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call408;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call408;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call408;
reg    ap_block_pp0_stage0_11001_ignoreCallOp509;
wire    call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_ready;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_0;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_1;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_2;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_3;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_4;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_5;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_6;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_7;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_8;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_9;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_10;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_11;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_12;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_13;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_14;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_15;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_16;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_17;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_18;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_19;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_20;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_21;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_22;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_23;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_24;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_25;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_26;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_27;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_28;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_29;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_30;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_31;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_32;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_33;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_34;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_35;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_36;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_37;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_38;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_39;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_40;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_41;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_42;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_43;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_44;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_45;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_46;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_47;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_48;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_49;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_50;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_51;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_52;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_53;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_54;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_55;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_56;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_57;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_58;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_59;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_60;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_61;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_62;
wire   [15:0] call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_63;
wire    call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_ready;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_0;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_1;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_2;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_3;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_4;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_5;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_6;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_7;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_8;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_9;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_10;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_11;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_12;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_13;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_14;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_15;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_16;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_17;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_18;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_19;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_20;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_21;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_22;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_23;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_24;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_25;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_26;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_27;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_28;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_29;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_30;
wire   [15:0] call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_31;
wire    call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_ready;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_0;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_1;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_2;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_3;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_4;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_5;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_6;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_7;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_8;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_9;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_10;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_11;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_12;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_13;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_14;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_15;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_16;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_17;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_18;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_19;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_20;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_21;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_22;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_23;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_24;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_25;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_26;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_27;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_28;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_29;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_30;
wire   [15:0] call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_31;
wire   [15:0] grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_0;
wire   [15:0] grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_1;
wire   [15:0] grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_2;
wire   [15:0] grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_3;
wire   [15:0] grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_4;
reg    grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_ce;
reg    ap_block_state1_pp0_stage0_iter0_ignore_call414;
wire    ap_block_state2_pp0_stage0_iter1_ignore_call414;
wire    ap_block_state3_pp0_stage0_iter2_ignore_call414;
wire    ap_block_state4_pp0_stage0_iter3_ignore_call414;
wire    ap_block_state5_pp0_stage0_iter4_ignore_call414;
wire    ap_block_state6_pp0_stage0_iter5_ignore_call414;
wire    ap_block_state7_pp0_stage0_iter6_ignore_call414;
wire    ap_block_state8_pp0_stage0_iter7_ignore_call414;
wire    ap_block_state9_pp0_stage0_iter8_ignore_call414;
wire    ap_block_state10_pp0_stage0_iter9_ignore_call414;
wire    ap_block_state11_pp0_stage0_iter10_ignore_call414;
wire    ap_block_state12_pp0_stage0_iter11_ignore_call414;
wire    ap_block_state13_pp0_stage0_iter12_ignore_call414;
wire    ap_block_state14_pp0_stage0_iter13_ignore_call414;
wire    ap_block_state15_pp0_stage0_iter14_ignore_call414;
wire    ap_block_state16_pp0_stage0_iter15_ignore_call414;
wire    ap_block_state17_pp0_stage0_iter16_ignore_call414;
wire    ap_block_state18_pp0_stage0_iter17_ignore_call414;
wire    ap_block_state19_pp0_stage0_iter18_ignore_call414;
wire    ap_block_state20_pp0_stage0_iter19_ignore_call414;
wire    ap_block_state21_pp0_stage0_iter20_ignore_call414;
wire    ap_block_state22_pp0_stage0_iter21_ignore_call414;
wire    ap_block_state23_pp0_stage0_iter22_ignore_call414;
wire    ap_block_state24_pp0_stage0_iter23_ignore_call414;
wire    ap_block_state25_pp0_stage0_iter24_ignore_call414;
wire    ap_block_state26_pp0_stage0_iter25_ignore_call414;
wire    ap_block_state27_pp0_stage0_iter26_ignore_call414;
wire    ap_block_state28_pp0_stage0_iter27_ignore_call414;
wire    ap_block_state29_pp0_stage0_iter28_ignore_call414;
wire    ap_block_state30_pp0_stage0_iter29_ignore_call414;
wire    ap_block_state31_pp0_stage0_iter30_ignore_call414;
wire    ap_block_state32_pp0_stage0_iter31_ignore_call414;
wire    ap_block_state33_pp0_stage0_iter32_ignore_call414;
wire    ap_block_state34_pp0_stage0_iter33_ignore_call414;
wire    ap_block_state35_pp0_stage0_iter34_ignore_call414;
wire    ap_block_state36_pp0_stage0_iter35_ignore_call414;
wire    ap_block_state37_pp0_stage0_iter36_ignore_call414;
wire    ap_block_state38_pp0_stage0_iter37_ignore_call414;
wire    ap_block_state39_pp0_stage0_iter38_ignore_call414;
wire    ap_block_state40_pp0_stage0_iter39_ignore_call414;
wire    ap_block_state41_pp0_stage0_iter40_ignore_call414;
wire    ap_block_state42_pp0_stage0_iter41_ignore_call414;
wire    ap_block_state43_pp0_stage0_iter42_ignore_call414;
wire    ap_block_state44_pp0_stage0_iter43_ignore_call414;
wire    ap_block_state45_pp0_stage0_iter44_ignore_call414;
wire    ap_block_state46_pp0_stage0_iter45_ignore_call414;
wire    ap_block_state47_pp0_stage0_iter46_ignore_call414;
wire    ap_block_state48_pp0_stage0_iter47_ignore_call414;
wire    ap_block_state49_pp0_stage0_iter48_ignore_call414;
wire    ap_block_state50_pp0_stage0_iter49_ignore_call414;
wire    ap_block_state51_pp0_stage0_iter50_ignore_call414;
wire    ap_block_state52_pp0_stage0_iter51_ignore_call414;
wire    ap_block_state53_pp0_stage0_iter52_ignore_call414;
wire    ap_block_state54_pp0_stage0_iter53_ignore_call414;
wire    ap_block_state55_pp0_stage0_iter54_ignore_call414;
wire    ap_block_state56_pp0_stage0_iter55_ignore_call414;
wire    ap_block_state57_pp0_stage0_iter56_ignore_call414;
wire    ap_block_state58_pp0_stage0_iter57_ignore_call414;
wire    ap_block_state59_pp0_stage0_iter58_ignore_call414;
wire    ap_block_state60_pp0_stage0_iter59_ignore_call414;
wire    ap_block_state61_pp0_stage0_iter60_ignore_call414;
wire    ap_block_state62_pp0_stage0_iter61_ignore_call414;
wire    ap_block_state63_pp0_stage0_iter62_ignore_call414;
wire    ap_block_state64_pp0_stage0_iter63_ignore_call414;
wire    ap_block_state65_pp0_stage0_iter64_ignore_call414;
wire    ap_block_state66_pp0_stage0_iter65_ignore_call414;
wire    ap_block_state67_pp0_stage0_iter66_ignore_call414;
wire    ap_block_state68_pp0_stage0_iter67_ignore_call414;
reg    ap_block_pp0_stage0_11001_ignoreCallOp523;
reg    ap_block_pp0_stage0_01001;
reg   [0:0] ap_NS_fsm;
reg    ap_idle_pp0_0to66;
reg    ap_reset_idle_pp0;
wire    ap_enable_pp0;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
#0 ap_enable_reg_pp0_iter23 = 1'b0;
#0 ap_enable_reg_pp0_iter24 = 1'b0;
#0 ap_enable_reg_pp0_iter25 = 1'b0;
#0 ap_enable_reg_pp0_iter26 = 1'b0;
#0 ap_enable_reg_pp0_iter27 = 1'b0;
#0 ap_enable_reg_pp0_iter28 = 1'b0;
#0 ap_enable_reg_pp0_iter29 = 1'b0;
#0 ap_enable_reg_pp0_iter30 = 1'b0;
#0 ap_enable_reg_pp0_iter31 = 1'b0;
#0 ap_enable_reg_pp0_iter32 = 1'b0;
#0 ap_enable_reg_pp0_iter33 = 1'b0;
#0 ap_enable_reg_pp0_iter34 = 1'b0;
#0 ap_enable_reg_pp0_iter35 = 1'b0;
#0 ap_enable_reg_pp0_iter36 = 1'b0;
#0 ap_enable_reg_pp0_iter37 = 1'b0;
#0 ap_enable_reg_pp0_iter38 = 1'b0;
#0 ap_enable_reg_pp0_iter39 = 1'b0;
#0 ap_enable_reg_pp0_iter40 = 1'b0;
#0 ap_enable_reg_pp0_iter41 = 1'b0;
#0 ap_enable_reg_pp0_iter42 = 1'b0;
#0 ap_enable_reg_pp0_iter43 = 1'b0;
#0 ap_enable_reg_pp0_iter44 = 1'b0;
#0 ap_enable_reg_pp0_iter45 = 1'b0;
#0 ap_enable_reg_pp0_iter46 = 1'b0;
#0 ap_enable_reg_pp0_iter47 = 1'b0;
#0 ap_enable_reg_pp0_iter48 = 1'b0;
#0 ap_enable_reg_pp0_iter49 = 1'b0;
#0 ap_enable_reg_pp0_iter50 = 1'b0;
#0 ap_enable_reg_pp0_iter51 = 1'b0;
#0 ap_enable_reg_pp0_iter52 = 1'b0;
#0 ap_enable_reg_pp0_iter53 = 1'b0;
#0 ap_enable_reg_pp0_iter54 = 1'b0;
#0 ap_enable_reg_pp0_iter55 = 1'b0;
#0 ap_enable_reg_pp0_iter56 = 1'b0;
#0 ap_enable_reg_pp0_iter57 = 1'b0;
#0 ap_enable_reg_pp0_iter58 = 1'b0;
#0 ap_enable_reg_pp0_iter59 = 1'b0;
#0 ap_enable_reg_pp0_iter60 = 1'b0;
#0 ap_enable_reg_pp0_iter61 = 1'b0;
#0 ap_enable_reg_pp0_iter62 = 1'b0;
#0 ap_enable_reg_pp0_iter63 = 1'b0;
#0 ap_enable_reg_pp0_iter64 = 1'b0;
#0 ap_enable_reg_pp0_iter65 = 1'b0;
#0 ap_enable_reg_pp0_iter66 = 1'b0;
#0 ap_enable_reg_pp0_iter67 = 1'b0;
#0 input1_V_preg = 256'd0;
#0 input1_V_ap_vld_preg = 1'b0;
end

dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer5_out_0_V_reg_2786),
    .data_1_V_read(layer5_out_1_V_reg_2791),
    .data_2_V_read(layer5_out_2_V_reg_2796),
    .data_3_V_read(layer5_out_3_V_reg_2801),
    .data_4_V_read(layer5_out_4_V_reg_2806),
    .data_5_V_read(layer5_out_5_V_reg_2811),
    .data_6_V_read(layer5_out_6_V_reg_2816),
    .data_7_V_read(layer5_out_7_V_reg_2821),
    .data_8_V_read(layer5_out_8_V_reg_2826),
    .data_9_V_read(layer5_out_9_V_reg_2831),
    .data_10_V_read(layer5_out_10_V_reg_2836),
    .data_11_V_read(layer5_out_11_V_reg_2841),
    .data_12_V_read(layer5_out_12_V_reg_2846),
    .data_13_V_read(layer5_out_13_V_reg_2851),
    .data_14_V_read(layer5_out_14_V_reg_2856),
    .data_15_V_read(layer5_out_15_V_reg_2861),
    .data_16_V_read(layer5_out_16_V_reg_2866),
    .data_17_V_read(layer5_out_17_V_reg_2871),
    .data_18_V_read(layer5_out_18_V_reg_2876),
    .data_19_V_read(layer5_out_19_V_reg_2881),
    .data_20_V_read(layer5_out_20_V_reg_2886),
    .data_21_V_read(layer5_out_21_V_reg_2891),
    .data_22_V_read(layer5_out_22_V_reg_2896),
    .data_23_V_read(layer5_out_23_V_reg_2901),
    .data_24_V_read(layer5_out_24_V_reg_2906),
    .data_25_V_read(layer5_out_25_V_reg_2911),
    .data_26_V_read(layer5_out_26_V_reg_2916),
    .data_27_V_read(layer5_out_27_V_reg_2921),
    .data_28_V_read(layer5_out_28_V_reg_2926),
    .data_29_V_read(layer5_out_29_V_reg_2931),
    .data_30_V_read(layer5_out_30_V_reg_2936),
    .data_31_V_read(layer5_out_31_V_reg_2941),
    .data_32_V_read(layer5_out_32_V_reg_2946),
    .data_33_V_read(layer5_out_33_V_reg_2951),
    .data_34_V_read(layer5_out_34_V_reg_2956),
    .data_35_V_read(layer5_out_35_V_reg_2961),
    .data_36_V_read(layer5_out_36_V_reg_2966),
    .data_37_V_read(layer5_out_37_V_reg_2971),
    .data_38_V_read(layer5_out_38_V_reg_2976),
    .data_39_V_read(layer5_out_39_V_reg_2981),
    .data_40_V_read(layer5_out_40_V_reg_2986),
    .data_41_V_read(layer5_out_41_V_reg_2991),
    .data_42_V_read(layer5_out_42_V_reg_2996),
    .data_43_V_read(layer5_out_43_V_reg_3001),
    .data_44_V_read(layer5_out_44_V_reg_3006),
    .data_45_V_read(layer5_out_45_V_reg_3011),
    .data_46_V_read(layer5_out_46_V_reg_3016),
    .data_47_V_read(layer5_out_47_V_reg_3021),
    .data_48_V_read(layer5_out_48_V_reg_3026),
    .data_49_V_read(layer5_out_49_V_reg_3031),
    .data_50_V_read(layer5_out_50_V_reg_3036),
    .data_51_V_read(layer5_out_51_V_reg_3041),
    .data_52_V_read(layer5_out_52_V_reg_3046),
    .data_53_V_read(layer5_out_53_V_reg_3051),
    .data_54_V_read(layer5_out_54_V_reg_3056),
    .data_55_V_read(layer5_out_55_V_reg_3061),
    .data_56_V_read(layer5_out_56_V_reg_3066),
    .data_57_V_read(layer5_out_57_V_reg_3071),
    .data_58_V_read(layer5_out_58_V_reg_3076),
    .data_59_V_read(layer5_out_59_V_reg_3081),
    .data_60_V_read(layer5_out_60_V_reg_3086),
    .data_61_V_read(layer5_out_61_V_reg_3091),
    .data_62_V_read(layer5_out_62_V_reg_3096),
    .data_63_V_read(layer5_out_63_V_reg_3101),
    .ap_return_0(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_0),
    .ap_return_1(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_1),
    .ap_return_2(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_2),
    .ap_return_3(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_3),
    .ap_return_4(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_4),
    .ap_return_5(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_5),
    .ap_return_6(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_6),
    .ap_return_7(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_7),
    .ap_return_8(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_8),
    .ap_return_9(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_9),
    .ap_return_10(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_10),
    .ap_return_11(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_11),
    .ap_return_12(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_12),
    .ap_return_13(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_13),
    .ap_return_14(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_14),
    .ap_return_15(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_15),
    .ap_return_16(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_16),
    .ap_return_17(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_17),
    .ap_return_18(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_18),
    .ap_return_19(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_19),
    .ap_return_20(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_20),
    .ap_return_21(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_21),
    .ap_return_22(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_22),
    .ap_return_23(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_23),
    .ap_return_24(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_24),
    .ap_return_25(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_25),
    .ap_return_26(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_26),
    .ap_return_27(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_27),
    .ap_return_28(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_28),
    .ap_return_29(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_29),
    .ap_return_30(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_30),
    .ap_return_31(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_31),
    .ap_ce(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_ce)
);

dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer9_out_0_V_reg_3426),
    .data_1_V_read(layer9_out_1_V_reg_3431),
    .data_2_V_read(layer9_out_2_V_reg_3436),
    .data_3_V_read(layer9_out_3_V_reg_3441),
    .data_4_V_read(layer9_out_4_V_reg_3446),
    .data_5_V_read(layer9_out_5_V_reg_3451),
    .data_6_V_read(layer9_out_6_V_reg_3456),
    .data_7_V_read(layer9_out_7_V_reg_3461),
    .data_8_V_read(layer9_out_8_V_reg_3466),
    .data_9_V_read(layer9_out_9_V_reg_3471),
    .data_10_V_read(layer9_out_10_V_reg_3476),
    .data_11_V_read(layer9_out_11_V_reg_3481),
    .data_12_V_read(layer9_out_12_V_reg_3486),
    .data_13_V_read(layer9_out_13_V_reg_3491),
    .data_14_V_read(layer9_out_14_V_reg_3496),
    .data_15_V_read(layer9_out_15_V_reg_3501),
    .data_16_V_read(layer9_out_16_V_reg_3506),
    .data_17_V_read(layer9_out_17_V_reg_3511),
    .data_18_V_read(layer9_out_18_V_reg_3516),
    .data_19_V_read(layer9_out_19_V_reg_3521),
    .data_20_V_read(layer9_out_20_V_reg_3526),
    .data_21_V_read(layer9_out_21_V_reg_3531),
    .data_22_V_read(layer9_out_22_V_reg_3536),
    .data_23_V_read(layer9_out_23_V_reg_3541),
    .data_24_V_read(layer9_out_24_V_reg_3546),
    .data_25_V_read(layer9_out_25_V_reg_3551),
    .data_26_V_read(layer9_out_26_V_reg_3556),
    .data_27_V_read(layer9_out_27_V_reg_3561),
    .data_28_V_read(layer9_out_28_V_reg_3566),
    .data_29_V_read(layer9_out_29_V_reg_3571),
    .data_30_V_read(layer9_out_30_V_reg_3576),
    .data_31_V_read(layer9_out_31_V_reg_3581),
    .ap_return_0(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_0),
    .ap_return_1(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_1),
    .ap_return_2(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_2),
    .ap_return_3(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_3),
    .ap_return_4(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_4),
    .ap_return_5(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_5),
    .ap_return_6(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_6),
    .ap_return_7(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_7),
    .ap_return_8(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_8),
    .ap_return_9(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_9),
    .ap_return_10(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_10),
    .ap_return_11(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_11),
    .ap_return_12(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_12),
    .ap_return_13(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_13),
    .ap_return_14(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_14),
    .ap_return_15(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_15),
    .ap_return_16(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_16),
    .ap_return_17(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_17),
    .ap_return_18(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_18),
    .ap_return_19(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_19),
    .ap_return_20(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_20),
    .ap_return_21(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_21),
    .ap_return_22(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_22),
    .ap_return_23(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_23),
    .ap_return_24(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_24),
    .ap_return_25(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_25),
    .ap_return_26(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_26),
    .ap_return_27(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_27),
    .ap_return_28(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_28),
    .ap_return_29(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_29),
    .ap_return_30(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_30),
    .ap_return_31(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_31),
    .ap_ce(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_ce)
);

dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_V_read(input1_V_in_sig),
    .ap_return_0(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_0),
    .ap_return_1(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_1),
    .ap_return_2(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_2),
    .ap_return_3(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_3),
    .ap_return_4(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_4),
    .ap_return_5(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_5),
    .ap_return_6(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_6),
    .ap_return_7(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_7),
    .ap_return_8(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_8),
    .ap_return_9(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_9),
    .ap_return_10(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_10),
    .ap_return_11(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_11),
    .ap_return_12(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_12),
    .ap_return_13(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_13),
    .ap_return_14(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_14),
    .ap_return_15(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_15),
    .ap_return_16(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_16),
    .ap_return_17(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_17),
    .ap_return_18(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_18),
    .ap_return_19(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_19),
    .ap_return_20(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_20),
    .ap_return_21(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_21),
    .ap_return_22(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_22),
    .ap_return_23(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_23),
    .ap_return_24(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_24),
    .ap_return_25(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_25),
    .ap_return_26(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_26),
    .ap_return_27(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_27),
    .ap_return_28(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_28),
    .ap_return_29(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_29),
    .ap_return_30(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_30),
    .ap_return_31(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_31),
    .ap_return_32(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_32),
    .ap_return_33(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_33),
    .ap_return_34(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_34),
    .ap_return_35(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_35),
    .ap_return_36(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_36),
    .ap_return_37(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_37),
    .ap_return_38(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_38),
    .ap_return_39(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_39),
    .ap_return_40(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_40),
    .ap_return_41(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_41),
    .ap_return_42(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_42),
    .ap_return_43(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_43),
    .ap_return_44(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_44),
    .ap_return_45(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_45),
    .ap_return_46(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_46),
    .ap_return_47(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_47),
    .ap_return_48(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_48),
    .ap_return_49(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_49),
    .ap_return_50(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_50),
    .ap_return_51(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_51),
    .ap_return_52(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_52),
    .ap_return_53(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_53),
    .ap_return_54(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_54),
    .ap_return_55(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_55),
    .ap_return_56(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_56),
    .ap_return_57(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_57),
    .ap_return_58(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_58),
    .ap_return_59(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_59),
    .ap_return_60(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_60),
    .ap_return_61(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_61),
    .ap_return_62(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_62),
    .ap_return_63(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_63),
    .ap_ce(grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_ce)
);

normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer2_out_0_V_reg_2146),
    .data_1_V_read(layer2_out_1_V_reg_2151),
    .data_2_V_read(layer2_out_2_V_reg_2156),
    .data_3_V_read(layer2_out_3_V_reg_2161),
    .data_4_V_read(layer2_out_4_V_reg_2166),
    .data_5_V_read(layer2_out_5_V_reg_2171),
    .data_6_V_read(layer2_out_6_V_reg_2176),
    .data_7_V_read(layer2_out_7_V_reg_2181),
    .data_8_V_read(layer2_out_8_V_reg_2186),
    .data_9_V_read(layer2_out_9_V_reg_2191),
    .data_10_V_read(layer2_out_10_V_reg_2196),
    .data_11_V_read(layer2_out_11_V_reg_2201),
    .data_12_V_read(layer2_out_12_V_reg_2206),
    .data_13_V_read(layer2_out_13_V_reg_2211),
    .data_14_V_read(layer2_out_14_V_reg_2216),
    .data_15_V_read(layer2_out_15_V_reg_2221),
    .data_16_V_read(layer2_out_16_V_reg_2226),
    .data_17_V_read(layer2_out_17_V_reg_2231),
    .data_18_V_read(layer2_out_18_V_reg_2236),
    .data_19_V_read(layer2_out_19_V_reg_2241),
    .data_20_V_read(layer2_out_20_V_reg_2246),
    .data_21_V_read(layer2_out_21_V_reg_2251),
    .data_22_V_read(layer2_out_22_V_reg_2256),
    .data_23_V_read(layer2_out_23_V_reg_2261),
    .data_24_V_read(layer2_out_24_V_reg_2266),
    .data_25_V_read(layer2_out_25_V_reg_2271),
    .data_26_V_read(layer2_out_26_V_reg_2276),
    .data_27_V_read(layer2_out_27_V_reg_2281),
    .data_28_V_read(layer2_out_28_V_reg_2286),
    .data_29_V_read(layer2_out_29_V_reg_2291),
    .data_30_V_read(layer2_out_30_V_reg_2296),
    .data_31_V_read(layer2_out_31_V_reg_2301),
    .data_32_V_read(layer2_out_32_V_reg_2306),
    .data_33_V_read(layer2_out_33_V_reg_2311),
    .data_34_V_read(layer2_out_34_V_reg_2316),
    .data_35_V_read(layer2_out_35_V_reg_2321),
    .data_36_V_read(layer2_out_36_V_reg_2326),
    .data_37_V_read(layer2_out_37_V_reg_2331),
    .data_38_V_read(layer2_out_38_V_reg_2336),
    .data_39_V_read(layer2_out_39_V_reg_2341),
    .data_40_V_read(layer2_out_40_V_reg_2346),
    .data_41_V_read(layer2_out_41_V_reg_2351),
    .data_42_V_read(layer2_out_42_V_reg_2356),
    .data_43_V_read(layer2_out_43_V_reg_2361),
    .data_44_V_read(layer2_out_44_V_reg_2366),
    .data_45_V_read(layer2_out_45_V_reg_2371),
    .data_46_V_read(layer2_out_46_V_reg_2376),
    .data_47_V_read(layer2_out_47_V_reg_2381),
    .data_48_V_read(layer2_out_48_V_reg_2386),
    .data_49_V_read(layer2_out_49_V_reg_2391),
    .data_50_V_read(layer2_out_50_V_reg_2396),
    .data_51_V_read(layer2_out_51_V_reg_2401),
    .data_52_V_read(layer2_out_52_V_reg_2406),
    .data_53_V_read(layer2_out_53_V_reg_2411),
    .data_54_V_read(layer2_out_54_V_reg_2416),
    .data_55_V_read(layer2_out_55_V_reg_2421),
    .data_56_V_read(layer2_out_56_V_reg_2426),
    .data_57_V_read(layer2_out_57_V_reg_2431),
    .data_58_V_read(layer2_out_58_V_reg_2436),
    .data_59_V_read(layer2_out_59_V_reg_2441),
    .data_60_V_read(layer2_out_60_V_reg_2446),
    .data_61_V_read(layer2_out_61_V_reg_2451),
    .data_62_V_read(layer2_out_62_V_reg_2456),
    .data_63_V_read(layer2_out_63_V_reg_2461),
    .ap_return_0(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_0),
    .ap_return_1(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_1),
    .ap_return_2(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_2),
    .ap_return_3(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_3),
    .ap_return_4(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_4),
    .ap_return_5(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_5),
    .ap_return_6(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_6),
    .ap_return_7(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_7),
    .ap_return_8(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_8),
    .ap_return_9(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_9),
    .ap_return_10(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_10),
    .ap_return_11(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_11),
    .ap_return_12(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_12),
    .ap_return_13(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_13),
    .ap_return_14(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_14),
    .ap_return_15(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_15),
    .ap_return_16(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_16),
    .ap_return_17(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_17),
    .ap_return_18(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_18),
    .ap_return_19(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_19),
    .ap_return_20(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_20),
    .ap_return_21(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_21),
    .ap_return_22(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_22),
    .ap_return_23(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_23),
    .ap_return_24(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_24),
    .ap_return_25(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_25),
    .ap_return_26(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_26),
    .ap_return_27(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_27),
    .ap_return_28(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_28),
    .ap_return_29(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_29),
    .ap_return_30(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_30),
    .ap_return_31(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_31),
    .ap_return_32(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_32),
    .ap_return_33(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_33),
    .ap_return_34(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_34),
    .ap_return_35(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_35),
    .ap_return_36(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_36),
    .ap_return_37(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_37),
    .ap_return_38(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_38),
    .ap_return_39(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_39),
    .ap_return_40(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_40),
    .ap_return_41(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_41),
    .ap_return_42(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_42),
    .ap_return_43(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_43),
    .ap_return_44(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_44),
    .ap_return_45(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_45),
    .ap_return_46(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_46),
    .ap_return_47(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_47),
    .ap_return_48(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_48),
    .ap_return_49(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_49),
    .ap_return_50(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_50),
    .ap_return_51(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_51),
    .ap_return_52(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_52),
    .ap_return_53(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_53),
    .ap_return_54(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_54),
    .ap_return_55(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_55),
    .ap_return_56(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_56),
    .ap_return_57(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_57),
    .ap_return_58(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_58),
    .ap_return_59(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_59),
    .ap_return_60(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_60),
    .ap_return_61(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_61),
    .ap_return_62(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_62),
    .ap_return_63(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_63),
    .ap_ce(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_ce)
);

normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer10_out_0_V_reg_3586),
    .data_1_V_read(layer10_out_1_V_reg_3591),
    .data_2_V_read(layer10_out_2_V_reg_3596),
    .data_3_V_read(layer10_out_3_V_reg_3601),
    .data_4_V_read(layer10_out_4_V_reg_3606),
    .data_5_V_read(layer10_out_5_V_reg_3611),
    .data_6_V_read(layer10_out_6_V_reg_3616),
    .data_7_V_read(layer10_out_7_V_reg_3621),
    .data_8_V_read(layer10_out_8_V_reg_3626),
    .data_9_V_read(layer10_out_9_V_reg_3631),
    .data_10_V_read(layer10_out_10_V_reg_3636),
    .data_11_V_read(layer10_out_11_V_reg_3641),
    .data_12_V_read(layer10_out_12_V_reg_3646),
    .data_13_V_read(layer10_out_13_V_reg_3651),
    .data_14_V_read(layer10_out_14_V_reg_3656),
    .data_15_V_read(layer10_out_15_V_reg_3661),
    .data_16_V_read(layer10_out_16_V_reg_3666),
    .data_17_V_read(layer10_out_17_V_reg_3671),
    .data_18_V_read(layer10_out_18_V_reg_3676),
    .data_19_V_read(layer10_out_19_V_reg_3681),
    .data_20_V_read(layer10_out_20_V_reg_3686),
    .data_21_V_read(layer10_out_21_V_reg_3691),
    .data_22_V_read(layer10_out_22_V_reg_3696),
    .data_23_V_read(layer10_out_23_V_reg_3701),
    .data_24_V_read(layer10_out_24_V_reg_3706),
    .data_25_V_read(layer10_out_25_V_reg_3711),
    .data_26_V_read(layer10_out_26_V_reg_3716),
    .data_27_V_read(layer10_out_27_V_reg_3721),
    .data_28_V_read(layer10_out_28_V_reg_3726),
    .data_29_V_read(layer10_out_29_V_reg_3731),
    .data_30_V_read(layer10_out_30_V_reg_3736),
    .data_31_V_read(layer10_out_31_V_reg_3741),
    .ap_return_0(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_0),
    .ap_return_1(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_1),
    .ap_return_2(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_2),
    .ap_return_3(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_3),
    .ap_return_4(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_4),
    .ap_return_5(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_5),
    .ap_return_6(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_6),
    .ap_return_7(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_7),
    .ap_return_8(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_8),
    .ap_return_9(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_9),
    .ap_return_10(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_10),
    .ap_return_11(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_11),
    .ap_return_12(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_12),
    .ap_return_13(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_13),
    .ap_return_14(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_14),
    .ap_return_15(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_15),
    .ap_return_16(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_16),
    .ap_return_17(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_17),
    .ap_return_18(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_18),
    .ap_return_19(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_19),
    .ap_return_20(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_20),
    .ap_return_21(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_21),
    .ap_return_22(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_22),
    .ap_return_23(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_23),
    .ap_return_24(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_24),
    .ap_return_25(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_25),
    .ap_return_26(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_26),
    .ap_return_27(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_27),
    .ap_return_28(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_28),
    .ap_return_29(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_29),
    .ap_return_30(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_30),
    .ap_return_31(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_31),
    .ap_ce(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_ce)
);

normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer6_out_0_V_reg_3106),
    .data_1_V_read(layer6_out_1_V_reg_3111),
    .data_2_V_read(layer6_out_2_V_reg_3116),
    .data_3_V_read(layer6_out_3_V_reg_3121),
    .data_4_V_read(layer6_out_4_V_reg_3126),
    .data_5_V_read(layer6_out_5_V_reg_3131),
    .data_6_V_read(layer6_out_6_V_reg_3136),
    .data_7_V_read(layer6_out_7_V_reg_3141),
    .data_8_V_read(layer6_out_8_V_reg_3146),
    .data_9_V_read(layer6_out_9_V_reg_3151),
    .data_10_V_read(layer6_out_10_V_reg_3156),
    .data_11_V_read(layer6_out_11_V_reg_3161),
    .data_12_V_read(layer6_out_12_V_reg_3166),
    .data_13_V_read(layer6_out_13_V_reg_3171),
    .data_14_V_read(layer6_out_14_V_reg_3176),
    .data_15_V_read(layer6_out_15_V_reg_3181),
    .data_16_V_read(layer6_out_16_V_reg_3186),
    .data_17_V_read(layer6_out_17_V_reg_3191),
    .data_18_V_read(layer6_out_18_V_reg_3196),
    .data_19_V_read(layer6_out_19_V_reg_3201),
    .data_20_V_read(layer6_out_20_V_reg_3206),
    .data_21_V_read(layer6_out_21_V_reg_3211),
    .data_22_V_read(layer6_out_22_V_reg_3216),
    .data_23_V_read(layer6_out_23_V_reg_3221),
    .data_24_V_read(layer6_out_24_V_reg_3226),
    .data_25_V_read(layer6_out_25_V_reg_3231),
    .data_26_V_read(layer6_out_26_V_reg_3236),
    .data_27_V_read(layer6_out_27_V_reg_3241),
    .data_28_V_read(layer6_out_28_V_reg_3246),
    .data_29_V_read(layer6_out_29_V_reg_3251),
    .data_30_V_read(layer6_out_30_V_reg_3256),
    .data_31_V_read(layer6_out_31_V_reg_3261),
    .ap_return_0(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_0),
    .ap_return_1(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_1),
    .ap_return_2(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_2),
    .ap_return_3(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_3),
    .ap_return_4(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_4),
    .ap_return_5(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_5),
    .ap_return_6(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_6),
    .ap_return_7(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_7),
    .ap_return_8(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_8),
    .ap_return_9(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_9),
    .ap_return_10(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_10),
    .ap_return_11(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_11),
    .ap_return_12(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_12),
    .ap_return_13(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_13),
    .ap_return_14(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_14),
    .ap_return_15(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_15),
    .ap_return_16(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_16),
    .ap_return_17(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_17),
    .ap_return_18(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_18),
    .ap_return_19(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_19),
    .ap_return_20(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_20),
    .ap_return_21(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_21),
    .ap_return_22(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_22),
    .ap_return_23(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_23),
    .ap_return_24(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_24),
    .ap_return_25(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_25),
    .ap_return_26(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_26),
    .ap_return_27(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_27),
    .ap_return_28(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_28),
    .ap_return_29(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_29),
    .ap_return_30(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_30),
    .ap_return_31(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_31),
    .ap_ce(grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_ce)
);

dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0 grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer13_out_0_V_reg_3906),
    .data_1_V_read(layer13_out_1_V_reg_3911),
    .data_2_V_read(layer13_out_2_V_reg_3916),
    .data_3_V_read(layer13_out_3_V_reg_3921),
    .data_4_V_read(layer13_out_4_V_reg_3926),
    .data_5_V_read(layer13_out_5_V_reg_3931),
    .data_6_V_read(layer13_out_6_V_reg_3936),
    .data_7_V_read(layer13_out_7_V_reg_3941),
    .data_8_V_read(layer13_out_8_V_reg_3946),
    .data_9_V_read(layer13_out_9_V_reg_3951),
    .data_10_V_read(layer13_out_10_V_reg_3956),
    .data_11_V_read(layer13_out_11_V_reg_3961),
    .data_12_V_read(layer13_out_12_V_reg_3966),
    .data_13_V_read(layer13_out_13_V_reg_3971),
    .data_14_V_read(layer13_out_14_V_reg_3976),
    .data_15_V_read(layer13_out_15_V_reg_3981),
    .data_16_V_read(layer13_out_16_V_reg_3986),
    .data_17_V_read(layer13_out_17_V_reg_3991),
    .data_18_V_read(layer13_out_18_V_reg_3996),
    .data_19_V_read(layer13_out_19_V_reg_4001),
    .data_20_V_read(layer13_out_20_V_reg_4006),
    .data_21_V_read(layer13_out_21_V_reg_4011),
    .data_22_V_read(layer13_out_22_V_reg_4016),
    .data_23_V_read(layer13_out_23_V_reg_4021),
    .data_24_V_read(layer13_out_24_V_reg_4026),
    .data_25_V_read(layer13_out_25_V_reg_4031),
    .data_26_V_read(layer13_out_26_V_reg_4036),
    .data_27_V_read(layer13_out_27_V_reg_4041),
    .data_28_V_read(layer13_out_28_V_reg_4046),
    .data_29_V_read(layer13_out_29_V_reg_4051),
    .data_30_V_read(layer13_out_30_V_reg_4056),
    .data_31_V_read(layer13_out_31_V_reg_4061),
    .ap_return_0(grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_0),
    .ap_return_1(grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_1),
    .ap_return_2(grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_2),
    .ap_return_3(grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_3),
    .ap_return_4(grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_4),
    .ap_ce(grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_ce)
);

relu_max_ap_fixed_ap_fixed_1_relu1_config5_s call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411(
    .ap_ready(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_ready),
    .data_0_V_read(layer4_out_0_V_reg_2466),
    .data_1_V_read(layer4_out_1_V_reg_2471),
    .data_2_V_read(layer4_out_2_V_reg_2476),
    .data_3_V_read(layer4_out_3_V_reg_2481),
    .data_4_V_read(layer4_out_4_V_reg_2486),
    .data_5_V_read(layer4_out_5_V_reg_2491),
    .data_6_V_read(layer4_out_6_V_reg_2496),
    .data_7_V_read(layer4_out_7_V_reg_2501),
    .data_8_V_read(layer4_out_8_V_reg_2506),
    .data_9_V_read(layer4_out_9_V_reg_2511),
    .data_10_V_read(layer4_out_10_V_reg_2516),
    .data_11_V_read(layer4_out_11_V_reg_2521),
    .data_12_V_read(layer4_out_12_V_reg_2526),
    .data_13_V_read(layer4_out_13_V_reg_2531),
    .data_14_V_read(layer4_out_14_V_reg_2536),
    .data_15_V_read(layer4_out_15_V_reg_2541),
    .data_16_V_read(layer4_out_16_V_reg_2546),
    .data_17_V_read(layer4_out_17_V_reg_2551),
    .data_18_V_read(layer4_out_18_V_reg_2556),
    .data_19_V_read(layer4_out_19_V_reg_2561),
    .data_20_V_read(layer4_out_20_V_reg_2566),
    .data_21_V_read(layer4_out_21_V_reg_2571),
    .data_22_V_read(layer4_out_22_V_reg_2576),
    .data_23_V_read(layer4_out_23_V_reg_2581),
    .data_24_V_read(layer4_out_24_V_reg_2586),
    .data_25_V_read(layer4_out_25_V_reg_2591),
    .data_26_V_read(layer4_out_26_V_reg_2596),
    .data_27_V_read(layer4_out_27_V_reg_2601),
    .data_28_V_read(layer4_out_28_V_reg_2606),
    .data_29_V_read(layer4_out_29_V_reg_2611),
    .data_30_V_read(layer4_out_30_V_reg_2616),
    .data_31_V_read(layer4_out_31_V_reg_2621),
    .data_32_V_read(layer4_out_32_V_reg_2626),
    .data_33_V_read(layer4_out_33_V_reg_2631),
    .data_34_V_read(layer4_out_34_V_reg_2636),
    .data_35_V_read(layer4_out_35_V_reg_2641),
    .data_36_V_read(layer4_out_36_V_reg_2646),
    .data_37_V_read(layer4_out_37_V_reg_2651),
    .data_38_V_read(layer4_out_38_V_reg_2656),
    .data_39_V_read(layer4_out_39_V_reg_2661),
    .data_40_V_read(layer4_out_40_V_reg_2666),
    .data_41_V_read(layer4_out_41_V_reg_2671),
    .data_42_V_read(layer4_out_42_V_reg_2676),
    .data_43_V_read(layer4_out_43_V_reg_2681),
    .data_44_V_read(layer4_out_44_V_reg_2686),
    .data_45_V_read(layer4_out_45_V_reg_2691),
    .data_46_V_read(layer4_out_46_V_reg_2696),
    .data_47_V_read(layer4_out_47_V_reg_2701),
    .data_48_V_read(layer4_out_48_V_reg_2706),
    .data_49_V_read(layer4_out_49_V_reg_2711),
    .data_50_V_read(layer4_out_50_V_reg_2716),
    .data_51_V_read(layer4_out_51_V_reg_2721),
    .data_52_V_read(layer4_out_52_V_reg_2726),
    .data_53_V_read(layer4_out_53_V_reg_2731),
    .data_54_V_read(layer4_out_54_V_reg_2736),
    .data_55_V_read(layer4_out_55_V_reg_2741),
    .data_56_V_read(layer4_out_56_V_reg_2746),
    .data_57_V_read(layer4_out_57_V_reg_2751),
    .data_58_V_read(layer4_out_58_V_reg_2756),
    .data_59_V_read(layer4_out_59_V_reg_2761),
    .data_60_V_read(layer4_out_60_V_reg_2766),
    .data_61_V_read(layer4_out_61_V_reg_2771),
    .data_62_V_read(layer4_out_62_V_reg_2776),
    .data_63_V_read(layer4_out_63_V_reg_2781),
    .ap_return_0(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_0),
    .ap_return_1(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_1),
    .ap_return_2(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_2),
    .ap_return_3(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_3),
    .ap_return_4(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_4),
    .ap_return_5(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_5),
    .ap_return_6(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_6),
    .ap_return_7(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_7),
    .ap_return_8(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_8),
    .ap_return_9(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_9),
    .ap_return_10(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_10),
    .ap_return_11(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_11),
    .ap_return_12(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_12),
    .ap_return_13(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_13),
    .ap_return_14(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_14),
    .ap_return_15(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_15),
    .ap_return_16(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_16),
    .ap_return_17(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_17),
    .ap_return_18(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_18),
    .ap_return_19(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_19),
    .ap_return_20(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_20),
    .ap_return_21(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_21),
    .ap_return_22(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_22),
    .ap_return_23(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_23),
    .ap_return_24(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_24),
    .ap_return_25(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_25),
    .ap_return_26(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_26),
    .ap_return_27(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_27),
    .ap_return_28(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_28),
    .ap_return_29(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_29),
    .ap_return_30(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_30),
    .ap_return_31(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_31),
    .ap_return_32(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_32),
    .ap_return_33(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_33),
    .ap_return_34(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_34),
    .ap_return_35(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_35),
    .ap_return_36(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_36),
    .ap_return_37(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_37),
    .ap_return_38(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_38),
    .ap_return_39(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_39),
    .ap_return_40(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_40),
    .ap_return_41(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_41),
    .ap_return_42(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_42),
    .ap_return_43(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_43),
    .ap_return_44(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_44),
    .ap_return_45(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_45),
    .ap_return_46(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_46),
    .ap_return_47(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_47),
    .ap_return_48(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_48),
    .ap_return_49(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_49),
    .ap_return_50(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_50),
    .ap_return_51(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_51),
    .ap_return_52(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_52),
    .ap_return_53(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_53),
    .ap_return_54(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_54),
    .ap_return_55(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_55),
    .ap_return_56(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_56),
    .ap_return_57(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_57),
    .ap_return_58(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_58),
    .ap_return_59(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_59),
    .ap_return_60(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_60),
    .ap_return_61(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_61),
    .ap_return_62(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_62),
    .ap_return_63(call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_63)
);

relu_max_ap_fixed_ap_fixed_1_relu1_config9_s call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479(
    .ap_ready(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_ready),
    .data_0_V_read(layer8_out_0_V_reg_3266),
    .data_1_V_read(layer8_out_1_V_reg_3271),
    .data_2_V_read(layer8_out_2_V_reg_3276),
    .data_3_V_read(layer8_out_3_V_reg_3281),
    .data_4_V_read(layer8_out_4_V_reg_3286),
    .data_5_V_read(layer8_out_5_V_reg_3291),
    .data_6_V_read(layer8_out_6_V_reg_3296),
    .data_7_V_read(layer8_out_7_V_reg_3301),
    .data_8_V_read(layer8_out_8_V_reg_3306),
    .data_9_V_read(layer8_out_9_V_reg_3311),
    .data_10_V_read(layer8_out_10_V_reg_3316),
    .data_11_V_read(layer8_out_11_V_reg_3321),
    .data_12_V_read(layer8_out_12_V_reg_3326),
    .data_13_V_read(layer8_out_13_V_reg_3331),
    .data_14_V_read(layer8_out_14_V_reg_3336),
    .data_15_V_read(layer8_out_15_V_reg_3341),
    .data_16_V_read(layer8_out_16_V_reg_3346),
    .data_17_V_read(layer8_out_17_V_reg_3351),
    .data_18_V_read(layer8_out_18_V_reg_3356),
    .data_19_V_read(layer8_out_19_V_reg_3361),
    .data_20_V_read(layer8_out_20_V_reg_3366),
    .data_21_V_read(layer8_out_21_V_reg_3371),
    .data_22_V_read(layer8_out_22_V_reg_3376),
    .data_23_V_read(layer8_out_23_V_reg_3381),
    .data_24_V_read(layer8_out_24_V_reg_3386),
    .data_25_V_read(layer8_out_25_V_reg_3391),
    .data_26_V_read(layer8_out_26_V_reg_3396),
    .data_27_V_read(layer8_out_27_V_reg_3401),
    .data_28_V_read(layer8_out_28_V_reg_3406),
    .data_29_V_read(layer8_out_29_V_reg_3411),
    .data_30_V_read(layer8_out_30_V_reg_3416),
    .data_31_V_read(layer8_out_31_V_reg_3421),
    .ap_return_0(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_0),
    .ap_return_1(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_1),
    .ap_return_2(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_2),
    .ap_return_3(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_3),
    .ap_return_4(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_4),
    .ap_return_5(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_5),
    .ap_return_6(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_6),
    .ap_return_7(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_7),
    .ap_return_8(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_8),
    .ap_return_9(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_9),
    .ap_return_10(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_10),
    .ap_return_11(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_11),
    .ap_return_12(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_12),
    .ap_return_13(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_13),
    .ap_return_14(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_14),
    .ap_return_15(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_15),
    .ap_return_16(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_16),
    .ap_return_17(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_17),
    .ap_return_18(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_18),
    .ap_return_19(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_19),
    .ap_return_20(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_20),
    .ap_return_21(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_21),
    .ap_return_22(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_22),
    .ap_return_23(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_23),
    .ap_return_24(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_24),
    .ap_return_25(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_25),
    .ap_return_26(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_26),
    .ap_return_27(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_27),
    .ap_return_28(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_28),
    .ap_return_29(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_29),
    .ap_return_30(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_30),
    .ap_return_31(call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_31)
);

relu_max_ap_fixed_ap_fixed_1_relu1_config13_s call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515(
    .ap_ready(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_ready),
    .data_0_V_read(layer12_out_0_V_reg_3746),
    .data_1_V_read(layer12_out_1_V_reg_3751),
    .data_2_V_read(layer12_out_2_V_reg_3756),
    .data_3_V_read(layer12_out_3_V_reg_3761),
    .data_4_V_read(layer12_out_4_V_reg_3766),
    .data_5_V_read(layer12_out_5_V_reg_3771),
    .data_6_V_read(layer12_out_6_V_reg_3776),
    .data_7_V_read(layer12_out_7_V_reg_3781),
    .data_8_V_read(layer12_out_8_V_reg_3786),
    .data_9_V_read(layer12_out_9_V_reg_3791),
    .data_10_V_read(layer12_out_10_V_reg_3796),
    .data_11_V_read(layer12_out_11_V_reg_3801),
    .data_12_V_read(layer12_out_12_V_reg_3806),
    .data_13_V_read(layer12_out_13_V_reg_3811),
    .data_14_V_read(layer12_out_14_V_reg_3816),
    .data_15_V_read(layer12_out_15_V_reg_3821),
    .data_16_V_read(layer12_out_16_V_reg_3826),
    .data_17_V_read(layer12_out_17_V_reg_3831),
    .data_18_V_read(layer12_out_18_V_reg_3836),
    .data_19_V_read(layer12_out_19_V_reg_3841),
    .data_20_V_read(layer12_out_20_V_reg_3846),
    .data_21_V_read(layer12_out_21_V_reg_3851),
    .data_22_V_read(layer12_out_22_V_reg_3856),
    .data_23_V_read(layer12_out_23_V_reg_3861),
    .data_24_V_read(layer12_out_24_V_reg_3866),
    .data_25_V_read(layer12_out_25_V_reg_3871),
    .data_26_V_read(layer12_out_26_V_reg_3876),
    .data_27_V_read(layer12_out_27_V_reg_3881),
    .data_28_V_read(layer12_out_28_V_reg_3886),
    .data_29_V_read(layer12_out_29_V_reg_3891),
    .data_30_V_read(layer12_out_30_V_reg_3896),
    .data_31_V_read(layer12_out_31_V_reg_3901),
    .ap_return_0(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_0),
    .ap_return_1(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_1),
    .ap_return_2(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_2),
    .ap_return_3(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_3),
    .ap_return_4(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_4),
    .ap_return_5(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_5),
    .ap_return_6(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_6),
    .ap_return_7(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_7),
    .ap_return_8(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_8),
    .ap_return_9(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_9),
    .ap_return_10(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_10),
    .ap_return_11(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_11),
    .ap_return_12(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_12),
    .ap_return_13(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_13),
    .ap_return_14(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_14),
    .ap_return_15(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_15),
    .ap_return_16(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_16),
    .ap_return_17(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_17),
    .ap_return_18(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_18),
    .ap_return_19(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_19),
    .ap_return_20(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_20),
    .ap_return_21(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_21),
    .ap_return_22(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_22),
    .ap_return_23(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_23),
    .ap_return_24(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_24),
    .ap_return_25(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_25),
    .ap_return_26(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_26),
    .ap_return_27(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_27),
    .ap_return_28(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_28),
    .ap_return_29(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_29),
    .ap_return_30(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_30),
    .ap_return_31(call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_31)
);

normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0 grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .data_0_V_read(layer14_out_0_V_reg_4066),
    .data_1_V_read(layer14_out_1_V_reg_4071),
    .data_2_V_read(layer14_out_2_V_reg_4076),
    .data_3_V_read(layer14_out_3_V_reg_4081),
    .data_4_V_read(layer14_out_4_V_reg_4086),
    .ap_return_0(grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_0),
    .ap_return_1(grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_1),
    .ap_return_2(grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_2),
    .ap_return_3(grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_3),
    .ap_return_4(grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_4),
    .ap_ce(grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_ce)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter23 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter24 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter25 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter26 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter27 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter28 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter29 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter30 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter30 <= ap_enable_reg_pp0_iter29;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter31 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter31 <= ap_enable_reg_pp0_iter30;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter32 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter32 <= ap_enable_reg_pp0_iter31;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter33 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter33 <= ap_enable_reg_pp0_iter32;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter34 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter34 <= ap_enable_reg_pp0_iter33;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter35 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter35 <= ap_enable_reg_pp0_iter34;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter36 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter36 <= ap_enable_reg_pp0_iter35;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter37 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter37 <= ap_enable_reg_pp0_iter36;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter38 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter38 <= ap_enable_reg_pp0_iter37;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter39 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter39 <= ap_enable_reg_pp0_iter38;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter40 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter40 <= ap_enable_reg_pp0_iter39;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter41 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter41 <= ap_enable_reg_pp0_iter40;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter42 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter42 <= ap_enable_reg_pp0_iter41;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter43 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter43 <= ap_enable_reg_pp0_iter42;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter44 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter44 <= ap_enable_reg_pp0_iter43;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter45 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter45 <= ap_enable_reg_pp0_iter44;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter46 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter46 <= ap_enable_reg_pp0_iter45;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter47 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter47 <= ap_enable_reg_pp0_iter46;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter48 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter48 <= ap_enable_reg_pp0_iter47;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter49 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter49 <= ap_enable_reg_pp0_iter48;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter50 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter50 <= ap_enable_reg_pp0_iter49;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter51 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter51 <= ap_enable_reg_pp0_iter50;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter52 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter52 <= ap_enable_reg_pp0_iter51;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter53 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter53 <= ap_enable_reg_pp0_iter52;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter54 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter54 <= ap_enable_reg_pp0_iter53;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter55 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter55 <= ap_enable_reg_pp0_iter54;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter56 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter56 <= ap_enable_reg_pp0_iter55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter57 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter57 <= ap_enable_reg_pp0_iter56;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter58 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter58 <= ap_enable_reg_pp0_iter57;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter59 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter59 <= ap_enable_reg_pp0_iter58;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter60 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter60 <= ap_enable_reg_pp0_iter59;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter61 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter61 <= ap_enable_reg_pp0_iter60;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter62 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter62 <= ap_enable_reg_pp0_iter61;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter63 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter63 <= ap_enable_reg_pp0_iter62;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter64 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter64 <= ap_enable_reg_pp0_iter63;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter65 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter65 <= ap_enable_reg_pp0_iter64;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter66 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter66 <= ap_enable_reg_pp0_iter65;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter67 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter67 <= ap_enable_reg_pp0_iter66;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        input1_V_ap_vld_preg <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            input1_V_ap_vld_preg <= 1'b0;
        end else if ((~((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0)) & (input1_V_ap_vld == 1'b1))) begin
            input1_V_ap_vld_preg <= input1_V_ap_vld;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        input1_V_preg <= 256'd0;
    end else begin
        if ((~((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0)) & (input1_V_ap_vld == 1'b1))) begin
            input1_V_preg <= input1_V;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        layer10_out_0_V_reg_3586 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_0;
        layer10_out_10_V_reg_3636 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_10;
        layer10_out_11_V_reg_3641 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_11;
        layer10_out_12_V_reg_3646 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_12;
        layer10_out_13_V_reg_3651 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_13;
        layer10_out_14_V_reg_3656 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_14;
        layer10_out_15_V_reg_3661 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_15;
        layer10_out_16_V_reg_3666 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_16;
        layer10_out_17_V_reg_3671 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_17;
        layer10_out_18_V_reg_3676 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_18;
        layer10_out_19_V_reg_3681 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_19;
        layer10_out_1_V_reg_3591 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_1;
        layer10_out_20_V_reg_3686 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_20;
        layer10_out_21_V_reg_3691 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_21;
        layer10_out_22_V_reg_3696 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_22;
        layer10_out_23_V_reg_3701 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_23;
        layer10_out_24_V_reg_3706 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_24;
        layer10_out_25_V_reg_3711 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_25;
        layer10_out_26_V_reg_3716 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_26;
        layer10_out_27_V_reg_3721 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_27;
        layer10_out_28_V_reg_3726 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_28;
        layer10_out_29_V_reg_3731 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_29;
        layer10_out_2_V_reg_3596 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_2;
        layer10_out_30_V_reg_3736 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_30;
        layer10_out_31_V_reg_3741 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_31;
        layer10_out_3_V_reg_3601 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_3;
        layer10_out_4_V_reg_3606 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_4;
        layer10_out_5_V_reg_3611 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_5;
        layer10_out_6_V_reg_3616 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_6;
        layer10_out_7_V_reg_3621 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_7;
        layer10_out_8_V_reg_3626 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_8;
        layer10_out_9_V_reg_3631 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_return_9;
        layer12_out_0_V_reg_3746 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_0;
        layer12_out_10_V_reg_3796 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_10;
        layer12_out_11_V_reg_3801 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_11;
        layer12_out_12_V_reg_3806 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_12;
        layer12_out_13_V_reg_3811 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_13;
        layer12_out_14_V_reg_3816 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_14;
        layer12_out_15_V_reg_3821 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_15;
        layer12_out_16_V_reg_3826 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_16;
        layer12_out_17_V_reg_3831 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_17;
        layer12_out_18_V_reg_3836 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_18;
        layer12_out_19_V_reg_3841 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_19;
        layer12_out_1_V_reg_3751 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_1;
        layer12_out_20_V_reg_3846 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_20;
        layer12_out_21_V_reg_3851 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_21;
        layer12_out_22_V_reg_3856 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_22;
        layer12_out_23_V_reg_3861 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_23;
        layer12_out_24_V_reg_3866 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_24;
        layer12_out_25_V_reg_3871 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_25;
        layer12_out_26_V_reg_3876 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_26;
        layer12_out_27_V_reg_3881 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_27;
        layer12_out_28_V_reg_3886 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_28;
        layer12_out_29_V_reg_3891 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_29;
        layer12_out_2_V_reg_3756 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_2;
        layer12_out_30_V_reg_3896 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_30;
        layer12_out_31_V_reg_3901 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_31;
        layer12_out_3_V_reg_3761 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_3;
        layer12_out_4_V_reg_3766 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_4;
        layer12_out_5_V_reg_3771 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_5;
        layer12_out_6_V_reg_3776 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_6;
        layer12_out_7_V_reg_3781 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_7;
        layer12_out_8_V_reg_3786 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_8;
        layer12_out_9_V_reg_3791 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_return_9;
        layer13_out_0_V_reg_3906 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_0;
        layer13_out_10_V_reg_3956 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_10;
        layer13_out_11_V_reg_3961 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_11;
        layer13_out_12_V_reg_3966 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_12;
        layer13_out_13_V_reg_3971 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_13;
        layer13_out_14_V_reg_3976 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_14;
        layer13_out_15_V_reg_3981 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_15;
        layer13_out_16_V_reg_3986 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_16;
        layer13_out_17_V_reg_3991 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_17;
        layer13_out_18_V_reg_3996 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_18;
        layer13_out_19_V_reg_4001 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_19;
        layer13_out_1_V_reg_3911 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_1;
        layer13_out_20_V_reg_4006 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_20;
        layer13_out_21_V_reg_4011 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_21;
        layer13_out_22_V_reg_4016 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_22;
        layer13_out_23_V_reg_4021 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_23;
        layer13_out_24_V_reg_4026 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_24;
        layer13_out_25_V_reg_4031 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_25;
        layer13_out_26_V_reg_4036 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_26;
        layer13_out_27_V_reg_4041 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_27;
        layer13_out_28_V_reg_4046 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_28;
        layer13_out_29_V_reg_4051 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_29;
        layer13_out_2_V_reg_3916 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_2;
        layer13_out_30_V_reg_4056 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_30;
        layer13_out_31_V_reg_4061 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_31;
        layer13_out_3_V_reg_3921 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_3;
        layer13_out_4_V_reg_3926 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_4;
        layer13_out_5_V_reg_3931 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_5;
        layer13_out_6_V_reg_3936 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_6;
        layer13_out_7_V_reg_3941 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_7;
        layer13_out_8_V_reg_3946 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_8;
        layer13_out_9_V_reg_3951 <= call_ret_i2_relu_max_ap_fixed_ap_fixed_1_relu1_config13_s_fu_515_ap_return_9;
        layer14_out_0_V_reg_4066 <= grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_0;
        layer14_out_1_V_reg_4071 <= grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_1;
        layer14_out_2_V_reg_4076 <= grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_2;
        layer14_out_3_V_reg_4081 <= grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_3;
        layer14_out_4_V_reg_4086 <= grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_return_4;
        layer2_out_0_V_reg_2146 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_0;
        layer2_out_10_V_reg_2196 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_10;
        layer2_out_11_V_reg_2201 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_11;
        layer2_out_12_V_reg_2206 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_12;
        layer2_out_13_V_reg_2211 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_13;
        layer2_out_14_V_reg_2216 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_14;
        layer2_out_15_V_reg_2221 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_15;
        layer2_out_16_V_reg_2226 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_16;
        layer2_out_17_V_reg_2231 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_17;
        layer2_out_18_V_reg_2236 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_18;
        layer2_out_19_V_reg_2241 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_19;
        layer2_out_1_V_reg_2151 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_1;
        layer2_out_20_V_reg_2246 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_20;
        layer2_out_21_V_reg_2251 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_21;
        layer2_out_22_V_reg_2256 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_22;
        layer2_out_23_V_reg_2261 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_23;
        layer2_out_24_V_reg_2266 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_24;
        layer2_out_25_V_reg_2271 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_25;
        layer2_out_26_V_reg_2276 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_26;
        layer2_out_27_V_reg_2281 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_27;
        layer2_out_28_V_reg_2286 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_28;
        layer2_out_29_V_reg_2291 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_29;
        layer2_out_2_V_reg_2156 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_2;
        layer2_out_30_V_reg_2296 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_30;
        layer2_out_31_V_reg_2301 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_31;
        layer2_out_32_V_reg_2306 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_32;
        layer2_out_33_V_reg_2311 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_33;
        layer2_out_34_V_reg_2316 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_34;
        layer2_out_35_V_reg_2321 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_35;
        layer2_out_36_V_reg_2326 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_36;
        layer2_out_37_V_reg_2331 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_37;
        layer2_out_38_V_reg_2336 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_38;
        layer2_out_39_V_reg_2341 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_39;
        layer2_out_3_V_reg_2161 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_3;
        layer2_out_40_V_reg_2346 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_40;
        layer2_out_41_V_reg_2351 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_41;
        layer2_out_42_V_reg_2356 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_42;
        layer2_out_43_V_reg_2361 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_43;
        layer2_out_44_V_reg_2366 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_44;
        layer2_out_45_V_reg_2371 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_45;
        layer2_out_46_V_reg_2376 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_46;
        layer2_out_47_V_reg_2381 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_47;
        layer2_out_48_V_reg_2386 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_48;
        layer2_out_49_V_reg_2391 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_49;
        layer2_out_4_V_reg_2166 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_4;
        layer2_out_50_V_reg_2396 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_50;
        layer2_out_51_V_reg_2401 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_51;
        layer2_out_52_V_reg_2406 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_52;
        layer2_out_53_V_reg_2411 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_53;
        layer2_out_54_V_reg_2416 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_54;
        layer2_out_55_V_reg_2421 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_55;
        layer2_out_56_V_reg_2426 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_56;
        layer2_out_57_V_reg_2431 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_57;
        layer2_out_58_V_reg_2436 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_58;
        layer2_out_59_V_reg_2441 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_59;
        layer2_out_5_V_reg_2171 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_5;
        layer2_out_60_V_reg_2446 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_60;
        layer2_out_61_V_reg_2451 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_61;
        layer2_out_62_V_reg_2456 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_62;
        layer2_out_63_V_reg_2461 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_63;
        layer2_out_6_V_reg_2176 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_6;
        layer2_out_7_V_reg_2181 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_7;
        layer2_out_8_V_reg_2186 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_8;
        layer2_out_9_V_reg_2191 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_return_9;
        layer4_out_0_V_reg_2466 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_0;
        layer4_out_10_V_reg_2516 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_10;
        layer4_out_11_V_reg_2521 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_11;
        layer4_out_12_V_reg_2526 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_12;
        layer4_out_13_V_reg_2531 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_13;
        layer4_out_14_V_reg_2536 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_14;
        layer4_out_15_V_reg_2541 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_15;
        layer4_out_16_V_reg_2546 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_16;
        layer4_out_17_V_reg_2551 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_17;
        layer4_out_18_V_reg_2556 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_18;
        layer4_out_19_V_reg_2561 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_19;
        layer4_out_1_V_reg_2471 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_1;
        layer4_out_20_V_reg_2566 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_20;
        layer4_out_21_V_reg_2571 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_21;
        layer4_out_22_V_reg_2576 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_22;
        layer4_out_23_V_reg_2581 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_23;
        layer4_out_24_V_reg_2586 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_24;
        layer4_out_25_V_reg_2591 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_25;
        layer4_out_26_V_reg_2596 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_26;
        layer4_out_27_V_reg_2601 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_27;
        layer4_out_28_V_reg_2606 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_28;
        layer4_out_29_V_reg_2611 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_29;
        layer4_out_2_V_reg_2476 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_2;
        layer4_out_30_V_reg_2616 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_30;
        layer4_out_31_V_reg_2621 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_31;
        layer4_out_32_V_reg_2626 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_32;
        layer4_out_33_V_reg_2631 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_33;
        layer4_out_34_V_reg_2636 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_34;
        layer4_out_35_V_reg_2641 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_35;
        layer4_out_36_V_reg_2646 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_36;
        layer4_out_37_V_reg_2651 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_37;
        layer4_out_38_V_reg_2656 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_38;
        layer4_out_39_V_reg_2661 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_39;
        layer4_out_3_V_reg_2481 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_3;
        layer4_out_40_V_reg_2666 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_40;
        layer4_out_41_V_reg_2671 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_41;
        layer4_out_42_V_reg_2676 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_42;
        layer4_out_43_V_reg_2681 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_43;
        layer4_out_44_V_reg_2686 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_44;
        layer4_out_45_V_reg_2691 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_45;
        layer4_out_46_V_reg_2696 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_46;
        layer4_out_47_V_reg_2701 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_47;
        layer4_out_48_V_reg_2706 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_48;
        layer4_out_49_V_reg_2711 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_49;
        layer4_out_4_V_reg_2486 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_4;
        layer4_out_50_V_reg_2716 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_50;
        layer4_out_51_V_reg_2721 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_51;
        layer4_out_52_V_reg_2726 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_52;
        layer4_out_53_V_reg_2731 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_53;
        layer4_out_54_V_reg_2736 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_54;
        layer4_out_55_V_reg_2741 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_55;
        layer4_out_56_V_reg_2746 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_56;
        layer4_out_57_V_reg_2751 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_57;
        layer4_out_58_V_reg_2756 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_58;
        layer4_out_59_V_reg_2761 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_59;
        layer4_out_5_V_reg_2491 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_5;
        layer4_out_60_V_reg_2766 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_60;
        layer4_out_61_V_reg_2771 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_61;
        layer4_out_62_V_reg_2776 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_62;
        layer4_out_63_V_reg_2781 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_63;
        layer4_out_6_V_reg_2496 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_6;
        layer4_out_7_V_reg_2501 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_7;
        layer4_out_8_V_reg_2506 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_8;
        layer4_out_9_V_reg_2511 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_return_9;
        layer5_out_0_V_reg_2786 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_0;
        layer5_out_10_V_reg_2836 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_10;
        layer5_out_11_V_reg_2841 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_11;
        layer5_out_12_V_reg_2846 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_12;
        layer5_out_13_V_reg_2851 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_13;
        layer5_out_14_V_reg_2856 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_14;
        layer5_out_15_V_reg_2861 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_15;
        layer5_out_16_V_reg_2866 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_16;
        layer5_out_17_V_reg_2871 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_17;
        layer5_out_18_V_reg_2876 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_18;
        layer5_out_19_V_reg_2881 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_19;
        layer5_out_1_V_reg_2791 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_1;
        layer5_out_20_V_reg_2886 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_20;
        layer5_out_21_V_reg_2891 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_21;
        layer5_out_22_V_reg_2896 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_22;
        layer5_out_23_V_reg_2901 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_23;
        layer5_out_24_V_reg_2906 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_24;
        layer5_out_25_V_reg_2911 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_25;
        layer5_out_26_V_reg_2916 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_26;
        layer5_out_27_V_reg_2921 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_27;
        layer5_out_28_V_reg_2926 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_28;
        layer5_out_29_V_reg_2931 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_29;
        layer5_out_2_V_reg_2796 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_2;
        layer5_out_30_V_reg_2936 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_30;
        layer5_out_31_V_reg_2941 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_31;
        layer5_out_32_V_reg_2946 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_32;
        layer5_out_33_V_reg_2951 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_33;
        layer5_out_34_V_reg_2956 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_34;
        layer5_out_35_V_reg_2961 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_35;
        layer5_out_36_V_reg_2966 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_36;
        layer5_out_37_V_reg_2971 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_37;
        layer5_out_38_V_reg_2976 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_38;
        layer5_out_39_V_reg_2981 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_39;
        layer5_out_3_V_reg_2801 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_3;
        layer5_out_40_V_reg_2986 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_40;
        layer5_out_41_V_reg_2991 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_41;
        layer5_out_42_V_reg_2996 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_42;
        layer5_out_43_V_reg_3001 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_43;
        layer5_out_44_V_reg_3006 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_44;
        layer5_out_45_V_reg_3011 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_45;
        layer5_out_46_V_reg_3016 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_46;
        layer5_out_47_V_reg_3021 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_47;
        layer5_out_48_V_reg_3026 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_48;
        layer5_out_49_V_reg_3031 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_49;
        layer5_out_4_V_reg_2806 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_4;
        layer5_out_50_V_reg_3036 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_50;
        layer5_out_51_V_reg_3041 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_51;
        layer5_out_52_V_reg_3046 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_52;
        layer5_out_53_V_reg_3051 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_53;
        layer5_out_54_V_reg_3056 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_54;
        layer5_out_55_V_reg_3061 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_55;
        layer5_out_56_V_reg_3066 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_56;
        layer5_out_57_V_reg_3071 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_57;
        layer5_out_58_V_reg_3076 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_58;
        layer5_out_59_V_reg_3081 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_59;
        layer5_out_5_V_reg_2811 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_5;
        layer5_out_60_V_reg_3086 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_60;
        layer5_out_61_V_reg_3091 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_61;
        layer5_out_62_V_reg_3096 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_62;
        layer5_out_63_V_reg_3101 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_63;
        layer5_out_6_V_reg_2816 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_6;
        layer5_out_7_V_reg_2821 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_7;
        layer5_out_8_V_reg_2826 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_8;
        layer5_out_9_V_reg_2831 <= call_ret_i_relu_max_ap_fixed_ap_fixed_1_relu1_config5_s_fu_411_ap_return_9;
        layer6_out_0_V_reg_3106 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_0;
        layer6_out_10_V_reg_3156 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_10;
        layer6_out_11_V_reg_3161 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_11;
        layer6_out_12_V_reg_3166 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_12;
        layer6_out_13_V_reg_3171 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_13;
        layer6_out_14_V_reg_3176 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_14;
        layer6_out_15_V_reg_3181 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_15;
        layer6_out_16_V_reg_3186 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_16;
        layer6_out_17_V_reg_3191 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_17;
        layer6_out_18_V_reg_3196 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_18;
        layer6_out_19_V_reg_3201 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_19;
        layer6_out_1_V_reg_3111 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_1;
        layer6_out_20_V_reg_3206 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_20;
        layer6_out_21_V_reg_3211 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_21;
        layer6_out_22_V_reg_3216 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_22;
        layer6_out_23_V_reg_3221 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_23;
        layer6_out_24_V_reg_3226 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_24;
        layer6_out_25_V_reg_3231 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_25;
        layer6_out_26_V_reg_3236 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_26;
        layer6_out_27_V_reg_3241 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_27;
        layer6_out_28_V_reg_3246 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_28;
        layer6_out_29_V_reg_3251 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_29;
        layer6_out_2_V_reg_3116 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_2;
        layer6_out_30_V_reg_3256 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_30;
        layer6_out_31_V_reg_3261 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_31;
        layer6_out_3_V_reg_3121 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_3;
        layer6_out_4_V_reg_3126 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_4;
        layer6_out_5_V_reg_3131 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_5;
        layer6_out_6_V_reg_3136 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_6;
        layer6_out_7_V_reg_3141 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_7;
        layer6_out_8_V_reg_3146 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_8;
        layer6_out_9_V_reg_3151 <= grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_return_9;
        layer8_out_0_V_reg_3266 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_0;
        layer8_out_10_V_reg_3316 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_10;
        layer8_out_11_V_reg_3321 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_11;
        layer8_out_12_V_reg_3326 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_12;
        layer8_out_13_V_reg_3331 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_13;
        layer8_out_14_V_reg_3336 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_14;
        layer8_out_15_V_reg_3341 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_15;
        layer8_out_16_V_reg_3346 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_16;
        layer8_out_17_V_reg_3351 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_17;
        layer8_out_18_V_reg_3356 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_18;
        layer8_out_19_V_reg_3361 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_19;
        layer8_out_1_V_reg_3271 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_1;
        layer8_out_20_V_reg_3366 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_20;
        layer8_out_21_V_reg_3371 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_21;
        layer8_out_22_V_reg_3376 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_22;
        layer8_out_23_V_reg_3381 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_23;
        layer8_out_24_V_reg_3386 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_24;
        layer8_out_25_V_reg_3391 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_25;
        layer8_out_26_V_reg_3396 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_26;
        layer8_out_27_V_reg_3401 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_27;
        layer8_out_28_V_reg_3406 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_28;
        layer8_out_29_V_reg_3411 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_29;
        layer8_out_2_V_reg_3276 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_2;
        layer8_out_30_V_reg_3416 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_30;
        layer8_out_31_V_reg_3421 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_31;
        layer8_out_3_V_reg_3281 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_3;
        layer8_out_4_V_reg_3286 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_4;
        layer8_out_5_V_reg_3291 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_5;
        layer8_out_6_V_reg_3296 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_6;
        layer8_out_7_V_reg_3301 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_7;
        layer8_out_8_V_reg_3306 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_8;
        layer8_out_9_V_reg_3311 <= grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_return_9;
        layer9_out_0_V_reg_3426 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_0;
        layer9_out_10_V_reg_3476 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_10;
        layer9_out_11_V_reg_3481 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_11;
        layer9_out_12_V_reg_3486 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_12;
        layer9_out_13_V_reg_3491 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_13;
        layer9_out_14_V_reg_3496 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_14;
        layer9_out_15_V_reg_3501 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_15;
        layer9_out_16_V_reg_3506 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_16;
        layer9_out_17_V_reg_3511 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_17;
        layer9_out_18_V_reg_3516 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_18;
        layer9_out_19_V_reg_3521 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_19;
        layer9_out_1_V_reg_3431 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_1;
        layer9_out_20_V_reg_3526 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_20;
        layer9_out_21_V_reg_3531 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_21;
        layer9_out_22_V_reg_3536 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_22;
        layer9_out_23_V_reg_3541 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_23;
        layer9_out_24_V_reg_3546 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_24;
        layer9_out_25_V_reg_3551 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_25;
        layer9_out_26_V_reg_3556 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_26;
        layer9_out_27_V_reg_3561 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_27;
        layer9_out_28_V_reg_3566 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_28;
        layer9_out_29_V_reg_3571 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_29;
        layer9_out_2_V_reg_3436 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_2;
        layer9_out_30_V_reg_3576 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_30;
        layer9_out_31_V_reg_3581 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_31;
        layer9_out_3_V_reg_3441 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_3;
        layer9_out_4_V_reg_3446 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_4;
        layer9_out_5_V_reg_3451 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_5;
        layer9_out_6_V_reg_3456 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_6;
        layer9_out_7_V_reg_3461 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_7;
        layer9_out_8_V_reg_3466 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_8;
        layer9_out_9_V_reg_3471 <= call_ret_i1_relu_max_ap_fixed_ap_fixed_1_relu1_config9_s_fu_479_ap_return_9;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter67 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter66 == 1'b0) & (ap_enable_reg_pp0_iter65 == 1'b0) & (ap_enable_reg_pp0_iter64 == 1'b0) & (ap_enable_reg_pp0_iter63 == 1'b0) & (ap_enable_reg_pp0_iter62 == 1'b0) & (ap_enable_reg_pp0_iter61 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter60 == 1'b0) & (ap_enable_reg_pp0_iter59 == 1'b0) & (ap_enable_reg_pp0_iter58 == 1'b0) & (ap_enable_reg_pp0_iter57 == 1'b0) & (ap_enable_reg_pp0_iter56 == 1'b0) & (ap_enable_reg_pp0_iter55 == 1'b0) & (ap_enable_reg_pp0_iter54 == 1'b0) & (ap_enable_reg_pp0_iter53 == 1'b0) & (ap_enable_reg_pp0_iter52 == 1'b0) & (ap_enable_reg_pp0_iter51 == 1'b0) & (ap_enable_reg_pp0_iter50 == 1'b0) & (ap_enable_reg_pp0_iter49 == 1'b0) & (ap_enable_reg_pp0_iter48 == 1'b0) & (ap_enable_reg_pp0_iter47 == 1'b0) & (ap_enable_reg_pp0_iter46 == 1'b0) & (ap_enable_reg_pp0_iter45 == 1'b0) & (ap_enable_reg_pp0_iter44 == 1'b0) & (ap_enable_reg_pp0_iter43 == 1'b0) & (ap_enable_reg_pp0_iter42 == 1'b0) & (ap_enable_reg_pp0_iter41 == 1'b0) & (ap_enable_reg_pp0_iter40 == 1'b0) & (ap_enable_reg_pp0_iter39 == 1'b0) & (ap_enable_reg_pp0_iter38 == 1'b0) & (ap_enable_reg_pp0_iter37 == 1'b0) & (ap_enable_reg_pp0_iter36 == 1'b0) & (ap_enable_reg_pp0_iter35 == 1'b0) & (ap_enable_reg_pp0_iter34 == 1'b0) & (ap_enable_reg_pp0_iter33 == 1'b0) & (ap_enable_reg_pp0_iter32 == 1'b0) & (ap_enable_reg_pp0_iter31 == 1'b0) & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter66 == 1'b0) & (ap_enable_reg_pp0_iter65 == 1'b0) & (ap_enable_reg_pp0_iter64 == 1'b0) & (ap_enable_reg_pp0_iter63 == 1'b0) & (ap_enable_reg_pp0_iter62 == 1'b0) & (ap_enable_reg_pp0_iter61 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter60 == 1'b0) & (ap_enable_reg_pp0_iter59 == 1'b0) & (ap_enable_reg_pp0_iter58 == 1'b0) & (ap_enable_reg_pp0_iter57 == 1'b0) & (ap_enable_reg_pp0_iter56 == 1'b0) & (ap_enable_reg_pp0_iter55 == 1'b0) & (ap_enable_reg_pp0_iter54 == 1'b0) & (ap_enable_reg_pp0_iter53 == 1'b0) & (ap_enable_reg_pp0_iter52 == 1'b0) & (ap_enable_reg_pp0_iter51 == 1'b0) & (ap_enable_reg_pp0_iter50 == 1'b0) & (ap_enable_reg_pp0_iter49 == 1'b0) & (ap_enable_reg_pp0_iter48 == 1'b0) & (ap_enable_reg_pp0_iter47 == 1'b0) & (ap_enable_reg_pp0_iter46 == 1'b0) & (ap_enable_reg_pp0_iter45 == 1'b0) & (ap_enable_reg_pp0_iter44 == 1'b0) & (ap_enable_reg_pp0_iter43 == 1'b0) & (ap_enable_reg_pp0_iter42 == 1'b0) & (ap_enable_reg_pp0_iter41 == 1'b0) & (ap_enable_reg_pp0_iter40 == 1'b0) & (ap_enable_reg_pp0_iter39 == 1'b0) & (ap_enable_reg_pp0_iter38 == 1'b0) & (ap_enable_reg_pp0_iter37 == 1'b0) & (ap_enable_reg_pp0_iter36 == 1'b0) & (ap_enable_reg_pp0_iter35 == 1'b0) & (ap_enable_reg_pp0_iter34 == 1'b0) & (ap_enable_reg_pp0_iter33 == 1'b0) & (ap_enable_reg_pp0_iter32 == 1'b0) & (ap_enable_reg_pp0_iter31 == 1'b0) & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
        ap_idle_pp0_0to66 = 1'b1;
    end else begin
        ap_idle_pp0_0to66 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (ap_idle_pp0_0to66 == 1'b1))) begin
        ap_reset_idle_pp0 = 1'b1;
    end else begin
        ap_reset_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        const_size_in_1_ap_vld = 1'b1;
    end else begin
        const_size_in_1_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        const_size_out_1_ap_vld = 1'b1;
    end else begin
        const_size_out_1_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp70) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_ce = 1'b1;
    end else begin
        grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_229_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp397) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_ce = 1'b1;
    end else begin
        grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_193_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp277) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_ce = 1'b1;
    end else begin
        grp_dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_125_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp509) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_ce = 1'b1;
    end else begin
        grp_dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0_fu_375_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp144) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_ce = 1'b1;
    end else begin
        grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1_fu_235_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp440) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_ce = 1'b1;
    end else begin
        grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2_fu_303_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp328) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_ce = 1'b1;
    end else begin
        grp_normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s_fu_339_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001_ignoreCallOp523) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_ce = 1'b1;
    end else begin
        grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_ce = 1'b0;
    end
end

always @ (*) begin
    if ((input1_V_ap_vld == 1'b1)) begin
        input1_V_ap_vld_in_sig = input1_V_ap_vld;
    end else begin
        input1_V_ap_vld_in_sig = input1_V_ap_vld_preg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        input1_V_blk_n = input1_V_ap_vld;
    end else begin
        input1_V_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((input1_V_ap_vld == 1'b1)) begin
        input1_V_in_sig = input1_V;
    end else begin
        input1_V_in_sig = input1_V_preg;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        layer16_out_0_V_ap_vld = 1'b1;
    end else begin
        layer16_out_0_V_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        layer16_out_1_V_ap_vld = 1'b1;
    end else begin
        layer16_out_1_V_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        layer16_out_2_V_ap_vld = 1'b1;
    end else begin
        layer16_out_2_V_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        layer16_out_3_V_ap_vld = 1'b1;
    end else begin
        layer16_out_3_V_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter67 == 1'b1))) begin
        layer16_out_4_V_ap_vld = 1'b1;
    end else begin
        layer16_out_4_V_ap_vld = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp144 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp277 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp328 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp397 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp440 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp509 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp523 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_11001_ignoreCallOp70 = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((ap_start == 1'b1) & ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0)));
end

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18_ignore_call80 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call15 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call210 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call243 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call309 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call342 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call408 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call414 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0_ignore_call80 = ((ap_start == 1'b0) | (input1_V_ap_vld_in_sig == 1'b0));
end

assign ap_block_state20_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage0_iter26_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage0_iter27_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage0_iter28_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage0_iter29_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage0_iter30_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage0_iter31_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage0_iter32_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage0_iter33_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage0_iter34_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage0_iter35_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage0_iter36_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage0_iter37_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage0_iter38_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage0_iter39_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage0_iter40_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage0_iter41_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage0_iter42_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage0_iter43_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage0_iter44_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage0_iter45_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage0_iter46_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage0_iter47_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage0_iter48_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage0_iter49_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage0_iter50_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage0_iter51_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage0_iter52_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage0_iter53_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage0_iter54_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage0_iter55_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage0_iter56_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage0_iter57_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage0_iter58_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage0_iter59_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage0_iter60_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage0_iter61_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage0_iter62_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage0_iter63_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage0_iter64_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage0_iter65_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage0_iter66_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage0_iter67_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call15 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call210 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call243 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call309 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call342 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call408 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call414 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8_ignore_call80 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start;

assign const_size_in_1 = 16'd16;

assign const_size_out_1 = 16'd5;

assign layer16_out_0_V = grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_0;

assign layer16_out_1_V = grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_1;

assign layer16_out_2_V = grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_2;

assign layer16_out_3_V = grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_3;

assign layer16_out_4_V = grp_normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0_fu_551_ap_return_4;

endmodule //myproject
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        data_32_V_read,
        data_33_V_read,
        data_34_V_read,
        data_35_V_read,
        data_36_V_read,
        data_37_V_read,
        data_38_V_read,
        data_39_V_read,
        data_40_V_read,
        data_41_V_read,
        data_42_V_read,
        data_43_V_read,
        data_44_V_read,
        data_45_V_read,
        data_46_V_read,
        data_47_V_read,
        data_48_V_read,
        data_49_V_read,
        data_50_V_read,
        data_51_V_read,
        data_52_V_read,
        data_53_V_read,
        data_54_V_read,
        data_55_V_read,
        data_56_V_read,
        data_57_V_read,
        data_58_V_read,
        data_59_V_read,
        data_60_V_read,
        data_61_V_read,
        data_62_V_read,
        data_63_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
input  [15:0] data_32_V_read;
input  [15:0] data_33_V_read;
input  [15:0] data_34_V_read;
input  [15:0] data_35_V_read;
input  [15:0] data_36_V_read;
input  [15:0] data_37_V_read;
input  [15:0] data_38_V_read;
input  [15:0] data_39_V_read;
input  [15:0] data_40_V_read;
input  [15:0] data_41_V_read;
input  [15:0] data_42_V_read;
input  [15:0] data_43_V_read;
input  [15:0] data_44_V_read;
input  [15:0] data_45_V_read;
input  [15:0] data_46_V_read;
input  [15:0] data_47_V_read;
input  [15:0] data_48_V_read;
input  [15:0] data_49_V_read;
input  [15:0] data_50_V_read;
input  [15:0] data_51_V_read;
input  [15:0] data_52_V_read;
input  [15:0] data_53_V_read;
input  [15:0] data_54_V_read;
input  [15:0] data_55_V_read;
input  [15:0] data_56_V_read;
input  [15:0] data_57_V_read;
input  [15:0] data_58_V_read;
input  [15:0] data_59_V_read;
input  [15:0] data_60_V_read;
input  [15:0] data_61_V_read;
input  [15:0] data_62_V_read;
input  [15:0] data_63_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
output  [15:0] ap_return_32;
output  [15:0] ap_return_33;
output  [15:0] ap_return_34;
output  [15:0] ap_return_35;
output  [15:0] ap_return_36;
output  [15:0] ap_return_37;
output  [15:0] ap_return_38;
output  [15:0] ap_return_39;
output  [15:0] ap_return_40;
output  [15:0] ap_return_41;
output  [15:0] ap_return_42;
output  [15:0] ap_return_43;
output  [15:0] ap_return_44;
output  [15:0] ap_return_45;
output  [15:0] ap_return_46;
output  [15:0] ap_return_47;
output  [15:0] ap_return_48;
output  [15:0] ap_return_49;
output  [15:0] ap_return_50;
output  [15:0] ap_return_51;
output  [15:0] ap_return_52;
output  [15:0] ap_return_53;
output  [15:0] ap_return_54;
output  [15:0] ap_return_55;
output  [15:0] ap_return_56;
output  [15:0] ap_return_57;
output  [15:0] ap_return_58;
output  [15:0] ap_return_59;
output  [15:0] ap_return_60;
output  [15:0] ap_return_61;
output  [15:0] ap_return_62;
output  [15:0] ap_return_63;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;
reg[15:0] ap_return_32;
reg[15:0] ap_return_33;
reg[15:0] ap_return_34;
reg[15:0] ap_return_35;
reg[15:0] ap_return_36;
reg[15:0] ap_return_37;
reg[15:0] ap_return_38;
reg[15:0] ap_return_39;
reg[15:0] ap_return_40;
reg[15:0] ap_return_41;
reg[15:0] ap_return_42;
reg[15:0] ap_return_43;
reg[15:0] ap_return_44;
reg[15:0] ap_return_45;
reg[15:0] ap_return_46;
reg[15:0] ap_return_47;
reg[15:0] ap_return_48;
reg[15:0] ap_return_49;
reg[15:0] ap_return_50;
reg[15:0] ap_return_51;
reg[15:0] ap_return_52;
reg[15:0] ap_return_53;
reg[15:0] ap_return_54;
reg[15:0] ap_return_55;
reg[15:0] ap_return_56;
reg[15:0] ap_return_57;
reg[15:0] ap_return_58;
reg[15:0] ap_return_59;
reg[15:0] ap_return_60;
reg[15:0] ap_return_61;
reg[15:0] ap_return_62;
reg[15:0] ap_return_63;

reg   [15:0] data_46_V_read_2_reg_18625;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_42_V_read_2_reg_18631;
reg   [15:0] data_39_V_read_2_reg_18637;
reg   [15:0] trunc_ln_reg_18948;
reg   [15:0] trunc_ln708_31_reg_18953;
reg   [15:0] trunc_ln708_32_reg_18958;
reg   [15:0] trunc_ln708_s_reg_18963;
reg   [15:0] trunc_ln708_33_reg_18968;
reg   [15:0] trunc_ln708_34_reg_18973;
reg   [15:0] trunc_ln708_35_reg_18978;
reg   [15:0] trunc_ln708_36_reg_18983;
reg   [15:0] trunc_ln708_37_reg_18988;
reg   [15:0] trunc_ln708_38_reg_18993;
reg   [15:0] trunc_ln708_39_reg_18998;
reg   [15:0] trunc_ln708_40_reg_19003;
reg   [15:0] trunc_ln708_41_reg_19008;
reg   [15:0] trunc_ln708_42_reg_19013;
reg   [15:0] trunc_ln708_43_reg_19018;
reg   [15:0] trunc_ln708_44_reg_19023;
reg   [15:0] trunc_ln708_45_reg_19028;
reg   [15:0] trunc_ln708_46_reg_19033;
reg   [15:0] trunc_ln708_47_reg_19038;
reg   [15:0] trunc_ln708_48_reg_19043;
reg   [15:0] trunc_ln708_49_reg_19048;
reg   [15:0] trunc_ln708_50_reg_19053;
reg   [15:0] trunc_ln708_51_reg_19058;
reg   [15:0] trunc_ln708_52_reg_19063;
reg   [15:0] trunc_ln708_53_reg_19068;
reg   [15:0] trunc_ln708_54_reg_19073;
reg   [15:0] trunc_ln708_55_reg_19078;
reg   [15:0] trunc_ln708_56_reg_19083;
reg   [15:0] trunc_ln708_57_reg_19088;
reg   [15:0] trunc_ln708_58_reg_19093;
reg   [15:0] trunc_ln708_59_reg_19098;
reg   [15:0] trunc_ln708_60_reg_19103;
reg   [15:0] trunc_ln708_61_reg_19108;
reg   [15:0] trunc_ln708_62_reg_19113;
reg   [15:0] trunc_ln708_63_reg_19118;
reg   [15:0] trunc_ln708_64_reg_19123;
reg   [15:0] trunc_ln708_65_reg_19128;
reg   [15:0] trunc_ln708_66_reg_19133;
reg   [15:0] trunc_ln708_67_reg_19138;
reg   [15:0] trunc_ln708_68_reg_19143;
reg   [15:0] trunc_ln708_69_reg_19148;
reg   [15:0] trunc_ln708_70_reg_19153;
reg   [15:0] trunc_ln708_71_reg_19158;
reg   [15:0] trunc_ln708_72_reg_19163;
reg   [15:0] trunc_ln708_73_reg_19168;
reg   [15:0] trunc_ln708_74_reg_19173;
reg   [15:0] trunc_ln708_75_reg_19178;
reg   [15:0] trunc_ln708_76_reg_19183;
reg   [15:0] trunc_ln708_77_reg_19188;
reg   [15:0] trunc_ln708_78_reg_19193;
reg   [15:0] trunc_ln708_79_reg_19198;
reg   [15:0] trunc_ln708_80_reg_19203;
reg   [15:0] trunc_ln708_81_reg_19208;
reg   [15:0] trunc_ln708_82_reg_19213;
reg   [15:0] trunc_ln708_83_reg_19218;
reg   [15:0] trunc_ln708_84_reg_19223;
reg   [15:0] trunc_ln708_85_reg_19228;
reg   [15:0] trunc_ln708_86_reg_19233;
reg   [15:0] trunc_ln708_87_reg_19238;
reg   [15:0] trunc_ln708_88_reg_19243;
reg   [15:0] trunc_ln708_89_reg_19248;
reg   [15:0] trunc_ln708_90_reg_19253;
reg   [15:0] trunc_ln708_91_reg_19258;
reg   [15:0] trunc_ln708_92_reg_19263;
wire   [11:0] grp_fu_804_p1;
wire    ap_block_pp0_stage0;
wire   [11:0] grp_fu_805_p1;
wire   [11:0] grp_fu_806_p1;
wire   [11:0] grp_fu_807_p1;
wire   [10:0] grp_fu_808_p1;
wire   [10:0] grp_fu_809_p1;
wire   [11:0] grp_fu_810_p1;
wire   [10:0] grp_fu_811_p1;
wire   [11:0] grp_fu_812_p1;
wire   [12:0] grp_fu_813_p1;
wire   [11:0] grp_fu_814_p1;
wire   [11:0] grp_fu_815_p1;
wire   [11:0] grp_fu_816_p1;
wire   [11:0] grp_fu_818_p1;
wire   [10:0] grp_fu_819_p1;
wire   [11:0] grp_fu_820_p1;
wire   [11:0] grp_fu_821_p1;
wire   [11:0] grp_fu_822_p1;
wire   [11:0] grp_fu_823_p1;
wire   [11:0] grp_fu_824_p1;
wire   [10:0] grp_fu_825_p1;
wire   [11:0] grp_fu_826_p1;
wire   [11:0] grp_fu_827_p1;
wire   [10:0] grp_fu_828_p1;
wire   [10:0] grp_fu_829_p1;
wire   [11:0] grp_fu_830_p1;
wire   [10:0] grp_fu_831_p1;
wire   [10:0] grp_fu_832_p1;
wire   [11:0] grp_fu_833_p1;
wire   [10:0] grp_fu_834_p1;
wire   [11:0] grp_fu_835_p1;
wire   [11:0] grp_fu_837_p1;
wire   [12:0] grp_fu_838_p1;
wire   [10:0] grp_fu_839_p1;
wire   [11:0] grp_fu_840_p1;
wire   [10:0] grp_fu_841_p1;
wire   [11:0] grp_fu_842_p1;
wire   [10:0] grp_fu_843_p1;
wire   [10:0] grp_fu_844_p1;
wire   [10:0] grp_fu_845_p1;
wire   [11:0] grp_fu_846_p1;
wire   [11:0] grp_fu_847_p1;
wire   [10:0] grp_fu_848_p1;
wire   [11:0] grp_fu_849_p1;
wire   [10:0] grp_fu_850_p1;
wire   [11:0] grp_fu_851_p1;
wire   [11:0] grp_fu_852_p1;
wire   [10:0] grp_fu_853_p1;
wire   [12:0] grp_fu_854_p1;
wire   [11:0] grp_fu_855_p1;
wire   [10:0] grp_fu_856_p1;
wire   [11:0] grp_fu_857_p1;
wire   [10:0] grp_fu_858_p1;
wire   [11:0] grp_fu_859_p1;
wire   [11:0] grp_fu_860_p1;
wire   [11:0] grp_fu_861_p1;
wire   [11:0] grp_fu_862_p1;
wire   [11:0] grp_fu_863_p1;
wire   [10:0] grp_fu_864_p1;
wire   [11:0] grp_fu_866_p1;
wire   [12:0] grp_fu_867_p1;
wire   [25:0] grp_fu_852_p2;
wire   [25:0] grp_fu_832_p2;
wire   [25:0] grp_fu_860_p2;
wire   [25:0] grp_fu_828_p2;
wire   [25:0] grp_fu_857_p2;
wire   [25:0] grp_fu_846_p2;
wire   [25:0] grp_fu_829_p2;
wire   [25:0] grp_fu_866_p2;
wire   [25:0] grp_fu_819_p2;
wire   [25:0] grp_fu_844_p2;
wire   [25:0] grp_fu_859_p2;
wire   [25:0] grp_fu_856_p2;
wire   [25:0] grp_fu_834_p2;
wire   [25:0] grp_fu_813_p2;
wire   [25:0] grp_fu_816_p2;
wire   [25:0] grp_fu_812_p2;
wire   [25:0] grp_fu_837_p2;
wire   [25:0] grp_fu_849_p2;
wire   [25:0] grp_fu_818_p2;
wire   [25:0] grp_fu_810_p2;
wire   [25:0] grp_fu_815_p2;
wire   [25:0] grp_fu_811_p2;
wire   [25:0] grp_fu_824_p2;
wire   [25:0] grp_fu_830_p2;
wire   [25:0] grp_fu_839_p2;
wire   [25:0] grp_fu_850_p2;
wire   [25:0] grp_fu_827_p2;
wire   [25:0] grp_fu_847_p2;
wire   [25:0] grp_fu_845_p2;
wire   [25:0] grp_fu_853_p2;
wire   [25:0] grp_fu_814_p2;
wire   [25:0] grp_fu_840_p2;
wire   [25:0] grp_fu_808_p2;
wire   [25:0] grp_fu_858_p2;
wire   [25:0] grp_fu_835_p2;
wire   [25:0] grp_fu_804_p2;
wire   [25:0] grp_fu_841_p2;
wire   [25:0] grp_fu_807_p2;
wire   [25:0] grp_fu_825_p2;
wire   [22:0] shl_ln1118_5_fu_17614_p3;
wire   [25:0] shl_ln_fu_17607_p3;
wire   [25:0] sext_ln1118_73_fu_17621_p1;
wire   [25:0] add_ln1118_fu_17625_p2;
wire   [25:0] grp_fu_867_p2;
wire   [25:0] grp_fu_822_p2;
wire   [25:0] sext_ln1118_76_fu_17661_p1;
wire   [25:0] shl_ln1118_6_fu_17664_p3;
wire   [25:0] add_ln1118_1_fu_17671_p2;
wire   [25:0] grp_fu_851_p2;
wire   [25:0] grp_fu_826_p2;
wire   [25:0] grp_fu_855_p2;
wire   [21:0] shl_ln1118_8_fu_17724_p3;
wire   [25:0] shl_ln1118_7_fu_17717_p3;
wire   [25:0] sext_ln1118_80_fu_17731_p1;
wire   [25:0] add_ln1118_2_fu_17735_p2;
wire   [25:0] grp_fu_838_p2;
wire   [25:0] grp_fu_861_p2;
wire   [25:0] grp_fu_843_p2;
wire   [25:0] grp_fu_862_p2;
wire   [25:0] grp_fu_863_p2;
wire   [25:0] grp_fu_823_p2;
wire   [25:0] grp_fu_848_p2;
wire   [25:0] grp_fu_854_p2;
wire   [25:0] grp_fu_821_p2;
wire   [25:0] grp_fu_831_p2;
wire   [25:0] grp_fu_864_p2;
wire   [25:0] grp_fu_809_p2;
wire   [25:0] grp_fu_842_p2;
wire   [25:0] grp_fu_805_p2;
wire   [25:0] grp_fu_833_p2;
wire   [25:0] grp_fu_806_p2;
wire   [25:0] grp_fu_820_p2;
wire   [15:0] add_ln703_fu_17921_p2;
wire   [15:0] add_ln703_36_fu_17926_p2;
wire   [15:0] add_ln703_37_fu_17931_p2;
wire   [15:0] add_ln703_38_fu_17936_p2;
wire   [15:0] add_ln703_39_fu_17941_p2;
wire   [15:0] add_ln703_40_fu_17946_p2;
wire   [15:0] add_ln703_41_fu_17951_p2;
wire   [15:0] add_ln703_42_fu_17956_p2;
wire   [15:0] add_ln703_43_fu_17961_p2;
wire   [15:0] add_ln703_44_fu_17966_p2;
wire   [15:0] add_ln703_45_fu_17971_p2;
wire   [15:0] add_ln703_46_fu_17976_p2;
wire   [15:0] add_ln703_47_fu_17981_p2;
wire   [15:0] add_ln703_48_fu_17986_p2;
wire   [15:0] add_ln703_49_fu_17991_p2;
wire   [15:0] add_ln703_50_fu_17996_p2;
wire   [15:0] add_ln703_51_fu_18001_p2;
wire   [15:0] add_ln703_52_fu_18006_p2;
wire   [15:0] add_ln703_53_fu_18011_p2;
wire   [15:0] add_ln703_54_fu_18016_p2;
wire   [15:0] add_ln703_55_fu_18021_p2;
wire   [15:0] add_ln703_56_fu_18026_p2;
wire   [15:0] add_ln703_57_fu_18031_p2;
wire   [15:0] add_ln703_58_fu_18036_p2;
wire   [15:0] add_ln703_59_fu_18041_p2;
wire   [15:0] add_ln703_60_fu_18046_p2;
wire   [15:0] add_ln703_61_fu_18051_p2;
wire   [15:0] add_ln703_62_fu_18056_p2;
wire   [15:0] add_ln703_63_fu_18061_p2;
wire   [15:0] add_ln703_64_fu_18066_p2;
wire   [15:0] add_ln703_65_fu_18071_p2;
wire   [15:0] add_ln703_66_fu_18076_p2;
wire   [15:0] add_ln703_67_fu_18081_p2;
wire   [15:0] add_ln703_68_fu_18086_p2;
wire   [15:0] add_ln703_69_fu_18091_p2;
wire   [15:0] add_ln703_70_fu_18096_p2;
wire   [15:0] add_ln703_71_fu_18101_p2;
wire   [15:0] add_ln703_72_fu_18106_p2;
wire   [15:0] add_ln703_73_fu_18111_p2;
wire   [15:0] add_ln703_74_fu_18116_p2;
wire   [15:0] add_ln703_75_fu_18121_p2;
wire   [15:0] add_ln703_76_fu_18126_p2;
wire   [15:0] add_ln703_77_fu_18131_p2;
wire   [15:0] add_ln703_78_fu_18136_p2;
wire   [15:0] add_ln703_79_fu_18141_p2;
wire   [15:0] add_ln703_80_fu_18146_p2;
wire   [15:0] add_ln703_81_fu_18151_p2;
wire   [15:0] add_ln703_82_fu_18156_p2;
wire   [15:0] add_ln703_83_fu_18161_p2;
wire   [15:0] add_ln703_84_fu_18166_p2;
wire   [15:0] add_ln703_85_fu_18171_p2;
wire   [15:0] add_ln703_86_fu_18176_p2;
wire   [15:0] add_ln703_87_fu_18181_p2;
wire   [15:0] add_ln703_88_fu_18186_p2;
wire   [15:0] add_ln703_89_fu_18191_p2;
wire   [15:0] add_ln703_90_fu_18196_p2;
wire   [15:0] add_ln703_91_fu_18201_p2;
wire   [15:0] add_ln703_92_fu_18206_p2;
wire   [15:0] add_ln703_93_fu_18211_p2;
wire   [15:0] add_ln703_94_fu_18216_p2;
wire   [15:0] add_ln703_95_fu_18221_p2;
wire   [15:0] add_ln703_96_fu_18226_p2;
wire   [15:0] add_ln703_97_fu_18231_p2;
wire   [15:0] add_ln703_98_fu_18236_p2;
reg    grp_fu_804_ce;
reg    grp_fu_805_ce;
reg    grp_fu_806_ce;
reg    grp_fu_807_ce;
reg    grp_fu_808_ce;
reg    grp_fu_809_ce;
reg    grp_fu_810_ce;
reg    grp_fu_811_ce;
reg    grp_fu_812_ce;
reg    grp_fu_813_ce;
reg    grp_fu_814_ce;
reg    grp_fu_815_ce;
reg    grp_fu_816_ce;
reg    grp_fu_818_ce;
reg    grp_fu_819_ce;
reg    grp_fu_820_ce;
reg    grp_fu_821_ce;
reg    grp_fu_822_ce;
reg    grp_fu_823_ce;
reg    grp_fu_824_ce;
reg    grp_fu_825_ce;
reg    grp_fu_826_ce;
reg    grp_fu_827_ce;
reg    grp_fu_828_ce;
reg    grp_fu_829_ce;
reg    grp_fu_830_ce;
reg    grp_fu_831_ce;
reg    grp_fu_832_ce;
reg    grp_fu_833_ce;
reg    grp_fu_834_ce;
reg    grp_fu_835_ce;
reg    grp_fu_837_ce;
reg    grp_fu_838_ce;
reg    grp_fu_839_ce;
reg    grp_fu_840_ce;
reg    grp_fu_841_ce;
reg    grp_fu_842_ce;
reg    grp_fu_843_ce;
reg    grp_fu_844_ce;
reg    grp_fu_845_ce;
reg    grp_fu_846_ce;
reg    grp_fu_847_ce;
reg    grp_fu_848_ce;
reg    grp_fu_849_ce;
reg    grp_fu_850_ce;
reg    grp_fu_851_ce;
reg    grp_fu_852_ce;
reg    grp_fu_853_ce;
reg    grp_fu_854_ce;
reg    grp_fu_855_ce;
reg    grp_fu_856_ce;
reg    grp_fu_857_ce;
reg    grp_fu_858_ce;
reg    grp_fu_859_ce;
reg    grp_fu_860_ce;
reg    grp_fu_861_ce;
reg    grp_fu_862_ce;
reg    grp_fu_863_ce;
reg    grp_fu_864_ce;
reg    grp_fu_866_ce;
reg    grp_fu_867_ce;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] data_32_V_read_int_reg;
reg   [15:0] data_33_V_read_int_reg;
reg   [15:0] data_34_V_read_int_reg;
reg   [15:0] data_35_V_read_int_reg;
reg   [15:0] data_36_V_read_int_reg;
reg   [15:0] data_37_V_read_int_reg;
reg   [15:0] data_38_V_read_int_reg;
reg   [15:0] data_39_V_read_int_reg;
reg   [15:0] data_40_V_read_int_reg;
reg   [15:0] data_41_V_read_int_reg;
reg   [15:0] data_42_V_read_int_reg;
reg   [15:0] data_43_V_read_int_reg;
reg   [15:0] data_44_V_read_int_reg;
reg   [15:0] data_45_V_read_int_reg;
reg   [15:0] data_46_V_read_int_reg;
reg   [15:0] data_47_V_read_int_reg;
reg   [15:0] data_48_V_read_int_reg;
reg   [15:0] data_49_V_read_int_reg;
reg   [15:0] data_50_V_read_int_reg;
reg   [15:0] data_51_V_read_int_reg;
reg   [15:0] data_52_V_read_int_reg;
reg   [15:0] data_53_V_read_int_reg;
reg   [15:0] data_54_V_read_int_reg;
reg   [15:0] data_55_V_read_int_reg;
reg   [15:0] data_56_V_read_int_reg;
reg   [15:0] data_57_V_read_int_reg;
reg   [15:0] data_58_V_read_int_reg;
reg   [15:0] data_59_V_read_int_reg;
reg   [15:0] data_60_V_read_int_reg;
reg   [15:0] data_61_V_read_int_reg;
reg   [15:0] data_62_V_read_int_reg;
reg   [15:0] data_63_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;
reg   [15:0] ap_return_32_int_reg;
reg   [15:0] ap_return_33_int_reg;
reg   [15:0] ap_return_34_int_reg;
reg   [15:0] ap_return_35_int_reg;
reg   [15:0] ap_return_36_int_reg;
reg   [15:0] ap_return_37_int_reg;
reg   [15:0] ap_return_38_int_reg;
reg   [15:0] ap_return_39_int_reg;
reg   [15:0] ap_return_40_int_reg;
reg   [15:0] ap_return_41_int_reg;
reg   [15:0] ap_return_42_int_reg;
reg   [15:0] ap_return_43_int_reg;
reg   [15:0] ap_return_44_int_reg;
reg   [15:0] ap_return_45_int_reg;
reg   [15:0] ap_return_46_int_reg;
reg   [15:0] ap_return_47_int_reg;
reg   [15:0] ap_return_48_int_reg;
reg   [15:0] ap_return_49_int_reg;
reg   [15:0] ap_return_50_int_reg;
reg   [15:0] ap_return_51_int_reg;
reg   [15:0] ap_return_52_int_reg;
reg   [15:0] ap_return_53_int_reg;
reg   [15:0] ap_return_54_int_reg;
reg   [15:0] ap_return_55_int_reg;
reg   [15:0] ap_return_56_int_reg;
reg   [15:0] ap_return_57_int_reg;
reg   [15:0] ap_return_58_int_reg;
reg   [15:0] ap_return_59_int_reg;
reg   [15:0] ap_return_60_int_reg;
reg   [15:0] ap_return_61_int_reg;
reg   [15:0] ap_return_62_int_reg;
reg   [15:0] ap_return_63_int_reg;

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U2(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_35_V_read_int_reg),
    .din1(grp_fu_804_p1),
    .ce(grp_fu_804_ce),
    .dout(grp_fu_804_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U3(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_60_V_read_int_reg),
    .din1(grp_fu_805_p1),
    .ce(grp_fu_805_ce),
    .dout(grp_fu_805_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U4(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_62_V_read_int_reg),
    .din1(grp_fu_806_p1),
    .ce(grp_fu_806_ce),
    .dout(grp_fu_806_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U5(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_37_V_read_int_reg),
    .din1(grp_fu_807_p1),
    .ce(grp_fu_807_ce),
    .dout(grp_fu_807_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U6(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_32_V_read_int_reg),
    .din1(grp_fu_808_p1),
    .ce(grp_fu_808_ce),
    .dout(grp_fu_808_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U7(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_58_V_read_int_reg),
    .din1(grp_fu_809_p1),
    .ce(grp_fu_809_ce),
    .dout(grp_fu_809_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U8(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_19_V_read_int_reg),
    .din1(grp_fu_810_p1),
    .ce(grp_fu_810_ce),
    .dout(grp_fu_810_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U9(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_21_V_read_int_reg),
    .din1(grp_fu_811_p1),
    .ce(grp_fu_811_ce),
    .dout(grp_fu_811_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U10(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_15_V_read_int_reg),
    .din1(grp_fu_812_p1),
    .ce(grp_fu_812_ce),
    .dout(grp_fu_812_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U11(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_13_V_read_int_reg),
    .din1(grp_fu_813_p1),
    .ce(grp_fu_813_ce),
    .dout(grp_fu_813_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U12(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_30_V_read_int_reg),
    .din1(grp_fu_814_p1),
    .ce(grp_fu_814_ce),
    .dout(grp_fu_814_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U13(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_20_V_read_int_reg),
    .din1(grp_fu_815_p1),
    .ce(grp_fu_815_ce),
    .dout(grp_fu_815_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U14(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_14_V_read_int_reg),
    .din1(grp_fu_816_p1),
    .ce(grp_fu_816_ce),
    .dout(grp_fu_816_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U15(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_18_V_read_int_reg),
    .din1(grp_fu_818_p1),
    .ce(grp_fu_818_ce),
    .dout(grp_fu_818_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U16(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_8_V_read_int_reg),
    .din1(grp_fu_819_p1),
    .ce(grp_fu_819_ce),
    .dout(grp_fu_819_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U17(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_63_V_read_int_reg),
    .din1(grp_fu_820_p1),
    .ce(grp_fu_820_ce),
    .dout(grp_fu_820_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U18(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_55_V_read_int_reg),
    .din1(grp_fu_821_p1),
    .ce(grp_fu_821_ce),
    .dout(grp_fu_821_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U19(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_41_V_read_int_reg),
    .din1(grp_fu_822_p1),
    .ce(grp_fu_822_ce),
    .dout(grp_fu_822_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U20(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_52_V_read_int_reg),
    .din1(grp_fu_823_p1),
    .ce(grp_fu_823_ce),
    .dout(grp_fu_823_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U21(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_22_V_read_int_reg),
    .din1(grp_fu_824_p1),
    .ce(grp_fu_824_ce),
    .dout(grp_fu_824_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U22(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_38_V_read_int_reg),
    .din1(grp_fu_825_p1),
    .ce(grp_fu_825_ce),
    .dout(grp_fu_825_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U23(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_44_V_read_int_reg),
    .din1(grp_fu_826_p1),
    .ce(grp_fu_826_ce),
    .dout(grp_fu_826_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U24(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_26_V_read_int_reg),
    .din1(grp_fu_827_p1),
    .ce(grp_fu_827_ce),
    .dout(grp_fu_827_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U25(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_3_V_read_int_reg),
    .din1(grp_fu_828_p1),
    .ce(grp_fu_828_ce),
    .dout(grp_fu_828_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U26(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_6_V_read_int_reg),
    .din1(grp_fu_829_p1),
    .ce(grp_fu_829_ce),
    .dout(grp_fu_829_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U27(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_23_V_read_int_reg),
    .din1(grp_fu_830_p1),
    .ce(grp_fu_830_ce),
    .dout(grp_fu_830_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U28(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_56_V_read_int_reg),
    .din1(grp_fu_831_p1),
    .ce(grp_fu_831_ce),
    .dout(grp_fu_831_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U29(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_1_V_read_int_reg),
    .din1(grp_fu_832_p1),
    .ce(grp_fu_832_ce),
    .dout(grp_fu_832_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U30(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_61_V_read_int_reg),
    .din1(grp_fu_833_p1),
    .ce(grp_fu_833_ce),
    .dout(grp_fu_833_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U31(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_12_V_read_int_reg),
    .din1(grp_fu_834_p1),
    .ce(grp_fu_834_ce),
    .dout(grp_fu_834_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U32(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_34_V_read_int_reg),
    .din1(grp_fu_835_p1),
    .ce(grp_fu_835_ce),
    .dout(grp_fu_835_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U33(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_16_V_read_int_reg),
    .din1(grp_fu_837_p1),
    .ce(grp_fu_837_ce),
    .dout(grp_fu_837_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U34(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_47_V_read_int_reg),
    .din1(grp_fu_838_p1),
    .ce(grp_fu_838_ce),
    .dout(grp_fu_838_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U35(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_24_V_read_int_reg),
    .din1(grp_fu_839_p1),
    .ce(grp_fu_839_ce),
    .dout(grp_fu_839_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U36(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_31_V_read_int_reg),
    .din1(grp_fu_840_p1),
    .ce(grp_fu_840_ce),
    .dout(grp_fu_840_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U37(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_36_V_read_int_reg),
    .din1(grp_fu_841_p1),
    .ce(grp_fu_841_ce),
    .dout(grp_fu_841_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U38(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_59_V_read_int_reg),
    .din1(grp_fu_842_p1),
    .ce(grp_fu_842_ce),
    .dout(grp_fu_842_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U39(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_49_V_read_int_reg),
    .din1(grp_fu_843_p1),
    .ce(grp_fu_843_ce),
    .dout(grp_fu_843_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U40(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_9_V_read_int_reg),
    .din1(grp_fu_844_p1),
    .ce(grp_fu_844_ce),
    .dout(grp_fu_844_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U41(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_28_V_read_int_reg),
    .din1(grp_fu_845_p1),
    .ce(grp_fu_845_ce),
    .dout(grp_fu_845_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U42(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_5_V_read_int_reg),
    .din1(grp_fu_846_p1),
    .ce(grp_fu_846_ce),
    .dout(grp_fu_846_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U43(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_27_V_read_int_reg),
    .din1(grp_fu_847_p1),
    .ce(grp_fu_847_ce),
    .dout(grp_fu_847_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U44(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_53_V_read_int_reg),
    .din1(grp_fu_848_p1),
    .ce(grp_fu_848_ce),
    .dout(grp_fu_848_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U45(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_17_V_read_int_reg),
    .din1(grp_fu_849_p1),
    .ce(grp_fu_849_ce),
    .dout(grp_fu_849_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U46(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_25_V_read_int_reg),
    .din1(grp_fu_850_p1),
    .ce(grp_fu_850_ce),
    .dout(grp_fu_850_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U47(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_43_V_read_int_reg),
    .din1(grp_fu_851_p1),
    .ce(grp_fu_851_ce),
    .dout(grp_fu_851_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U48(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_0_V_read_int_reg),
    .din1(grp_fu_852_p1),
    .ce(grp_fu_852_ce),
    .dout(grp_fu_852_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U49(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_29_V_read_int_reg),
    .din1(grp_fu_853_p1),
    .ce(grp_fu_853_ce),
    .dout(grp_fu_853_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U50(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_54_V_read_int_reg),
    .din1(grp_fu_854_p1),
    .ce(grp_fu_854_ce),
    .dout(grp_fu_854_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U51(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_45_V_read_int_reg),
    .din1(grp_fu_855_p1),
    .ce(grp_fu_855_ce),
    .dout(grp_fu_855_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U52(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_11_V_read_int_reg),
    .din1(grp_fu_856_p1),
    .ce(grp_fu_856_ce),
    .dout(grp_fu_856_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U53(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_4_V_read_int_reg),
    .din1(grp_fu_857_p1),
    .ce(grp_fu_857_ce),
    .dout(grp_fu_857_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U54(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_33_V_read_int_reg),
    .din1(grp_fu_858_p1),
    .ce(grp_fu_858_ce),
    .dout(grp_fu_858_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U55(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_10_V_read_int_reg),
    .din1(grp_fu_859_p1),
    .ce(grp_fu_859_ce),
    .dout(grp_fu_859_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U56(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_2_V_read_int_reg),
    .din1(grp_fu_860_p1),
    .ce(grp_fu_860_ce),
    .dout(grp_fu_860_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U57(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_48_V_read_int_reg),
    .din1(grp_fu_861_p1),
    .ce(grp_fu_861_ce),
    .dout(grp_fu_861_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U58(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_50_V_read_int_reg),
    .din1(grp_fu_862_p1),
    .ce(grp_fu_862_ce),
    .dout(grp_fu_862_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U59(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_51_V_read_int_reg),
    .din1(grp_fu_863_p1),
    .ce(grp_fu_863_ce),
    .dout(grp_fu_863_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U60(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_57_V_read_int_reg),
    .din1(grp_fu_864_p1),
    .ce(grp_fu_864_ce),
    .dout(grp_fu_864_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U61(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_7_V_read_int_reg),
    .din1(grp_fu_866_p1),
    .ce(grp_fu_866_ce),
    .dout(grp_fu_866_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U62(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_40_V_read_int_reg),
    .din1(grp_fu_867_p1),
    .ce(grp_fu_867_ce),
    .dout(grp_fu_867_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_fu_17921_p2;
        ap_return_10_int_reg <= add_ln703_45_fu_17971_p2;
        ap_return_11_int_reg <= add_ln703_46_fu_17976_p2;
        ap_return_12_int_reg <= add_ln703_47_fu_17981_p2;
        ap_return_13_int_reg <= add_ln703_48_fu_17986_p2;
        ap_return_14_int_reg <= add_ln703_49_fu_17991_p2;
        ap_return_15_int_reg <= add_ln703_50_fu_17996_p2;
        ap_return_16_int_reg <= add_ln703_51_fu_18001_p2;
        ap_return_17_int_reg <= add_ln703_52_fu_18006_p2;
        ap_return_18_int_reg <= add_ln703_53_fu_18011_p2;
        ap_return_19_int_reg <= add_ln703_54_fu_18016_p2;
        ap_return_1_int_reg <= add_ln703_36_fu_17926_p2;
        ap_return_20_int_reg <= add_ln703_55_fu_18021_p2;
        ap_return_21_int_reg <= add_ln703_56_fu_18026_p2;
        ap_return_22_int_reg <= add_ln703_57_fu_18031_p2;
        ap_return_23_int_reg <= add_ln703_58_fu_18036_p2;
        ap_return_24_int_reg <= add_ln703_59_fu_18041_p2;
        ap_return_25_int_reg <= add_ln703_60_fu_18046_p2;
        ap_return_26_int_reg <= add_ln703_61_fu_18051_p2;
        ap_return_27_int_reg <= add_ln703_62_fu_18056_p2;
        ap_return_28_int_reg <= add_ln703_63_fu_18061_p2;
        ap_return_29_int_reg <= add_ln703_64_fu_18066_p2;
        ap_return_2_int_reg <= add_ln703_37_fu_17931_p2;
        ap_return_30_int_reg <= add_ln703_65_fu_18071_p2;
        ap_return_31_int_reg <= add_ln703_66_fu_18076_p2;
        ap_return_32_int_reg <= add_ln703_67_fu_18081_p2;
        ap_return_33_int_reg <= add_ln703_68_fu_18086_p2;
        ap_return_34_int_reg <= add_ln703_69_fu_18091_p2;
        ap_return_35_int_reg <= add_ln703_70_fu_18096_p2;
        ap_return_36_int_reg <= add_ln703_71_fu_18101_p2;
        ap_return_37_int_reg <= add_ln703_72_fu_18106_p2;
        ap_return_38_int_reg <= add_ln703_73_fu_18111_p2;
        ap_return_39_int_reg <= add_ln703_74_fu_18116_p2;
        ap_return_3_int_reg <= add_ln703_38_fu_17936_p2;
        ap_return_40_int_reg <= add_ln703_75_fu_18121_p2;
        ap_return_41_int_reg <= add_ln703_76_fu_18126_p2;
        ap_return_42_int_reg <= add_ln703_77_fu_18131_p2;
        ap_return_43_int_reg <= add_ln703_78_fu_18136_p2;
        ap_return_44_int_reg <= add_ln703_79_fu_18141_p2;
        ap_return_45_int_reg <= add_ln703_80_fu_18146_p2;
        ap_return_46_int_reg <= add_ln703_81_fu_18151_p2;
        ap_return_47_int_reg <= add_ln703_82_fu_18156_p2;
        ap_return_48_int_reg <= add_ln703_83_fu_18161_p2;
        ap_return_49_int_reg <= add_ln703_84_fu_18166_p2;
        ap_return_4_int_reg <= add_ln703_39_fu_17941_p2;
        ap_return_50_int_reg <= add_ln703_85_fu_18171_p2;
        ap_return_51_int_reg <= add_ln703_86_fu_18176_p2;
        ap_return_52_int_reg <= add_ln703_87_fu_18181_p2;
        ap_return_53_int_reg <= add_ln703_88_fu_18186_p2;
        ap_return_54_int_reg <= add_ln703_89_fu_18191_p2;
        ap_return_55_int_reg <= add_ln703_90_fu_18196_p2;
        ap_return_56_int_reg <= add_ln703_91_fu_18201_p2;
        ap_return_57_int_reg <= add_ln703_92_fu_18206_p2;
        ap_return_58_int_reg <= add_ln703_93_fu_18211_p2;
        ap_return_59_int_reg <= add_ln703_94_fu_18216_p2;
        ap_return_5_int_reg <= add_ln703_40_fu_17946_p2;
        ap_return_60_int_reg <= add_ln703_95_fu_18221_p2;
        ap_return_61_int_reg <= add_ln703_96_fu_18226_p2;
        ap_return_62_int_reg <= add_ln703_97_fu_18231_p2;
        ap_return_63_int_reg <= add_ln703_98_fu_18236_p2;
        ap_return_6_int_reg <= add_ln703_41_fu_17951_p2;
        ap_return_7_int_reg <= add_ln703_42_fu_17956_p2;
        ap_return_8_int_reg <= add_ln703_43_fu_17961_p2;
        ap_return_9_int_reg <= add_ln703_44_fu_17966_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_32_V_read_int_reg <= data_32_V_read;
        data_33_V_read_int_reg <= data_33_V_read;
        data_34_V_read_int_reg <= data_34_V_read;
        data_35_V_read_int_reg <= data_35_V_read;
        data_36_V_read_int_reg <= data_36_V_read;
        data_37_V_read_int_reg <= data_37_V_read;
        data_38_V_read_int_reg <= data_38_V_read;
        data_39_V_read_int_reg <= data_39_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_40_V_read_int_reg <= data_40_V_read;
        data_41_V_read_int_reg <= data_41_V_read;
        data_42_V_read_int_reg <= data_42_V_read;
        data_43_V_read_int_reg <= data_43_V_read;
        data_44_V_read_int_reg <= data_44_V_read;
        data_45_V_read_int_reg <= data_45_V_read;
        data_46_V_read_int_reg <= data_46_V_read;
        data_47_V_read_int_reg <= data_47_V_read;
        data_48_V_read_int_reg <= data_48_V_read;
        data_49_V_read_int_reg <= data_49_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_50_V_read_int_reg <= data_50_V_read;
        data_51_V_read_int_reg <= data_51_V_read;
        data_52_V_read_int_reg <= data_52_V_read;
        data_53_V_read_int_reg <= data_53_V_read;
        data_54_V_read_int_reg <= data_54_V_read;
        data_55_V_read_int_reg <= data_55_V_read;
        data_56_V_read_int_reg <= data_56_V_read;
        data_57_V_read_int_reg <= data_57_V_read;
        data_58_V_read_int_reg <= data_58_V_read;
        data_59_V_read_int_reg <= data_59_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_60_V_read_int_reg <= data_60_V_read;
        data_61_V_read_int_reg <= data_61_V_read;
        data_62_V_read_int_reg <= data_62_V_read;
        data_63_V_read_int_reg <= data_63_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        data_39_V_read_2_reg_18637 <= data_39_V_read_int_reg;
        data_42_V_read_2_reg_18631 <= data_42_V_read_int_reg;
        data_46_V_read_2_reg_18625 <= data_46_V_read_int_reg;
        trunc_ln708_31_reg_18953 <= {{grp_fu_832_p2[25:10]}};
        trunc_ln708_32_reg_18958 <= {{grp_fu_860_p2[25:10]}};
        trunc_ln708_33_reg_18968 <= {{grp_fu_857_p2[25:10]}};
        trunc_ln708_34_reg_18973 <= {{grp_fu_846_p2[25:10]}};
        trunc_ln708_35_reg_18978 <= {{grp_fu_829_p2[25:10]}};
        trunc_ln708_36_reg_18983 <= {{grp_fu_866_p2[25:10]}};
        trunc_ln708_37_reg_18988 <= {{grp_fu_819_p2[25:10]}};
        trunc_ln708_38_reg_18993 <= {{grp_fu_844_p2[25:10]}};
        trunc_ln708_39_reg_18998 <= {{grp_fu_859_p2[25:10]}};
        trunc_ln708_40_reg_19003 <= {{grp_fu_856_p2[25:10]}};
        trunc_ln708_41_reg_19008 <= {{grp_fu_834_p2[25:10]}};
        trunc_ln708_42_reg_19013 <= {{grp_fu_813_p2[25:10]}};
        trunc_ln708_43_reg_19018 <= {{grp_fu_816_p2[25:10]}};
        trunc_ln708_44_reg_19023 <= {{grp_fu_812_p2[25:10]}};
        trunc_ln708_45_reg_19028 <= {{grp_fu_837_p2[25:10]}};
        trunc_ln708_46_reg_19033 <= {{grp_fu_849_p2[25:10]}};
        trunc_ln708_47_reg_19038 <= {{grp_fu_818_p2[25:10]}};
        trunc_ln708_48_reg_19043 <= {{grp_fu_810_p2[25:10]}};
        trunc_ln708_49_reg_19048 <= {{grp_fu_815_p2[25:10]}};
        trunc_ln708_50_reg_19053 <= {{grp_fu_811_p2[25:10]}};
        trunc_ln708_51_reg_19058 <= {{grp_fu_824_p2[25:10]}};
        trunc_ln708_52_reg_19063 <= {{grp_fu_830_p2[25:10]}};
        trunc_ln708_53_reg_19068 <= {{grp_fu_839_p2[25:10]}};
        trunc_ln708_54_reg_19073 <= {{grp_fu_850_p2[25:10]}};
        trunc_ln708_55_reg_19078 <= {{grp_fu_827_p2[25:10]}};
        trunc_ln708_56_reg_19083 <= {{grp_fu_847_p2[25:10]}};
        trunc_ln708_57_reg_19088 <= {{grp_fu_845_p2[25:10]}};
        trunc_ln708_58_reg_19093 <= {{grp_fu_853_p2[25:10]}};
        trunc_ln708_59_reg_19098 <= {{grp_fu_814_p2[25:10]}};
        trunc_ln708_60_reg_19103 <= {{grp_fu_840_p2[25:10]}};
        trunc_ln708_61_reg_19108 <= {{grp_fu_808_p2[25:10]}};
        trunc_ln708_62_reg_19113 <= {{grp_fu_858_p2[25:10]}};
        trunc_ln708_63_reg_19118 <= {{grp_fu_835_p2[25:10]}};
        trunc_ln708_64_reg_19123 <= {{grp_fu_804_p2[25:10]}};
        trunc_ln708_65_reg_19128 <= {{grp_fu_841_p2[25:10]}};
        trunc_ln708_66_reg_19133 <= {{grp_fu_807_p2[25:10]}};
        trunc_ln708_67_reg_19138 <= {{grp_fu_825_p2[25:10]}};
        trunc_ln708_68_reg_19143 <= {{add_ln1118_fu_17625_p2[25:10]}};
        trunc_ln708_69_reg_19148 <= {{grp_fu_867_p2[25:10]}};
        trunc_ln708_70_reg_19153 <= {{grp_fu_822_p2[25:10]}};
        trunc_ln708_71_reg_19158 <= {{add_ln1118_1_fu_17671_p2[25:10]}};
        trunc_ln708_72_reg_19163 <= {{grp_fu_851_p2[25:10]}};
        trunc_ln708_73_reg_19168 <= {{grp_fu_826_p2[25:10]}};
        trunc_ln708_74_reg_19173 <= {{grp_fu_855_p2[25:10]}};
        trunc_ln708_75_reg_19178 <= {{add_ln1118_2_fu_17735_p2[25:10]}};
        trunc_ln708_76_reg_19183 <= {{grp_fu_838_p2[25:10]}};
        trunc_ln708_77_reg_19188 <= {{grp_fu_861_p2[25:10]}};
        trunc_ln708_78_reg_19193 <= {{grp_fu_843_p2[25:10]}};
        trunc_ln708_79_reg_19198 <= {{grp_fu_862_p2[25:10]}};
        trunc_ln708_80_reg_19203 <= {{grp_fu_863_p2[25:10]}};
        trunc_ln708_81_reg_19208 <= {{grp_fu_823_p2[25:10]}};
        trunc_ln708_82_reg_19213 <= {{grp_fu_848_p2[25:10]}};
        trunc_ln708_83_reg_19218 <= {{grp_fu_854_p2[25:10]}};
        trunc_ln708_84_reg_19223 <= {{grp_fu_821_p2[25:10]}};
        trunc_ln708_85_reg_19228 <= {{grp_fu_831_p2[25:10]}};
        trunc_ln708_86_reg_19233 <= {{grp_fu_864_p2[25:10]}};
        trunc_ln708_87_reg_19238 <= {{grp_fu_809_p2[25:10]}};
        trunc_ln708_88_reg_19243 <= {{grp_fu_842_p2[25:10]}};
        trunc_ln708_89_reg_19248 <= {{grp_fu_805_p2[25:10]}};
        trunc_ln708_90_reg_19253 <= {{grp_fu_833_p2[25:10]}};
        trunc_ln708_91_reg_19258 <= {{grp_fu_806_p2[25:10]}};
        trunc_ln708_92_reg_19263 <= {{grp_fu_820_p2[25:10]}};
        trunc_ln708_s_reg_18963 <= {{grp_fu_828_p2[25:10]}};
        trunc_ln_reg_18948 <= {{grp_fu_852_p2[25:10]}};
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_fu_17921_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = add_ln703_36_fu_17926_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = add_ln703_45_fu_17971_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = add_ln703_46_fu_17976_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = add_ln703_47_fu_17981_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = add_ln703_48_fu_17986_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = add_ln703_49_fu_17991_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = add_ln703_50_fu_17996_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = add_ln703_51_fu_18001_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = add_ln703_52_fu_18006_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = add_ln703_53_fu_18011_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = add_ln703_54_fu_18016_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = add_ln703_37_fu_17931_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = add_ln703_55_fu_18021_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = add_ln703_56_fu_18026_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = add_ln703_57_fu_18031_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = add_ln703_58_fu_18036_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = add_ln703_59_fu_18041_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = add_ln703_60_fu_18046_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = add_ln703_61_fu_18051_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = add_ln703_62_fu_18056_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = add_ln703_63_fu_18061_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = add_ln703_64_fu_18066_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = add_ln703_38_fu_17936_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = add_ln703_65_fu_18071_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = add_ln703_66_fu_18076_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_32 = ap_return_32_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_32 = add_ln703_67_fu_18081_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_33 = ap_return_33_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_33 = add_ln703_68_fu_18086_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_34 = ap_return_34_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_34 = add_ln703_69_fu_18091_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_35 = ap_return_35_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_35 = add_ln703_70_fu_18096_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_36 = ap_return_36_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_36 = add_ln703_71_fu_18101_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_37 = ap_return_37_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_37 = add_ln703_72_fu_18106_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_38 = ap_return_38_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_38 = add_ln703_73_fu_18111_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_39 = ap_return_39_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_39 = add_ln703_74_fu_18116_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = add_ln703_39_fu_17941_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_40 = ap_return_40_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_40 = add_ln703_75_fu_18121_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_41 = ap_return_41_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_41 = add_ln703_76_fu_18126_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_42 = ap_return_42_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_42 = add_ln703_77_fu_18131_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_43 = ap_return_43_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_43 = add_ln703_78_fu_18136_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_44 = ap_return_44_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_44 = add_ln703_79_fu_18141_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_45 = ap_return_45_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_45 = add_ln703_80_fu_18146_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_46 = ap_return_46_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_46 = add_ln703_81_fu_18151_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_47 = ap_return_47_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_47 = add_ln703_82_fu_18156_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_48 = ap_return_48_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_48 = add_ln703_83_fu_18161_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_49 = ap_return_49_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_49 = add_ln703_84_fu_18166_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = add_ln703_40_fu_17946_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_50 = ap_return_50_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_50 = add_ln703_85_fu_18171_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_51 = ap_return_51_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_51 = add_ln703_86_fu_18176_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_52 = ap_return_52_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_52 = add_ln703_87_fu_18181_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_53 = ap_return_53_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_53 = add_ln703_88_fu_18186_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_54 = ap_return_54_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_54 = add_ln703_89_fu_18191_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_55 = ap_return_55_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_55 = add_ln703_90_fu_18196_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_56 = ap_return_56_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_56 = add_ln703_91_fu_18201_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_57 = ap_return_57_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_57 = add_ln703_92_fu_18206_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_58 = ap_return_58_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_58 = add_ln703_93_fu_18211_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_59 = ap_return_59_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_59 = add_ln703_94_fu_18216_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = add_ln703_41_fu_17951_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_60 = ap_return_60_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_60 = add_ln703_95_fu_18221_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_61 = ap_return_61_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_61 = add_ln703_96_fu_18226_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_62 = ap_return_62_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_62 = add_ln703_97_fu_18231_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_63 = ap_return_63_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_63 = add_ln703_98_fu_18236_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = add_ln703_42_fu_17956_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = add_ln703_43_fu_17961_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = add_ln703_44_fu_17966_p2;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_804_ce = 1'b1;
    end else begin
        grp_fu_804_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_805_ce = 1'b1;
    end else begin
        grp_fu_805_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_806_ce = 1'b1;
    end else begin
        grp_fu_806_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_807_ce = 1'b1;
    end else begin
        grp_fu_807_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_808_ce = 1'b1;
    end else begin
        grp_fu_808_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_809_ce = 1'b1;
    end else begin
        grp_fu_809_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_810_ce = 1'b1;
    end else begin
        grp_fu_810_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_811_ce = 1'b1;
    end else begin
        grp_fu_811_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_812_ce = 1'b1;
    end else begin
        grp_fu_812_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_813_ce = 1'b1;
    end else begin
        grp_fu_813_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_814_ce = 1'b1;
    end else begin
        grp_fu_814_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_815_ce = 1'b1;
    end else begin
        grp_fu_815_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_816_ce = 1'b1;
    end else begin
        grp_fu_816_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_818_ce = 1'b1;
    end else begin
        grp_fu_818_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_819_ce = 1'b1;
    end else begin
        grp_fu_819_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_820_ce = 1'b1;
    end else begin
        grp_fu_820_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_821_ce = 1'b1;
    end else begin
        grp_fu_821_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_822_ce = 1'b1;
    end else begin
        grp_fu_822_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_823_ce = 1'b1;
    end else begin
        grp_fu_823_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_824_ce = 1'b1;
    end else begin
        grp_fu_824_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_825_ce = 1'b1;
    end else begin
        grp_fu_825_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_826_ce = 1'b1;
    end else begin
        grp_fu_826_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_827_ce = 1'b1;
    end else begin
        grp_fu_827_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_828_ce = 1'b1;
    end else begin
        grp_fu_828_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_829_ce = 1'b1;
    end else begin
        grp_fu_829_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_830_ce = 1'b1;
    end else begin
        grp_fu_830_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_831_ce = 1'b1;
    end else begin
        grp_fu_831_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_832_ce = 1'b1;
    end else begin
        grp_fu_832_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_833_ce = 1'b1;
    end else begin
        grp_fu_833_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_834_ce = 1'b1;
    end else begin
        grp_fu_834_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_835_ce = 1'b1;
    end else begin
        grp_fu_835_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_837_ce = 1'b1;
    end else begin
        grp_fu_837_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_838_ce = 1'b1;
    end else begin
        grp_fu_838_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_839_ce = 1'b1;
    end else begin
        grp_fu_839_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_840_ce = 1'b1;
    end else begin
        grp_fu_840_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_841_ce = 1'b1;
    end else begin
        grp_fu_841_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_842_ce = 1'b1;
    end else begin
        grp_fu_842_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_843_ce = 1'b1;
    end else begin
        grp_fu_843_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_844_ce = 1'b1;
    end else begin
        grp_fu_844_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_845_ce = 1'b1;
    end else begin
        grp_fu_845_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_846_ce = 1'b1;
    end else begin
        grp_fu_846_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_847_ce = 1'b1;
    end else begin
        grp_fu_847_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_848_ce = 1'b1;
    end else begin
        grp_fu_848_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_849_ce = 1'b1;
    end else begin
        grp_fu_849_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_850_ce = 1'b1;
    end else begin
        grp_fu_850_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_851_ce = 1'b1;
    end else begin
        grp_fu_851_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_852_ce = 1'b1;
    end else begin
        grp_fu_852_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_853_ce = 1'b1;
    end else begin
        grp_fu_853_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_854_ce = 1'b1;
    end else begin
        grp_fu_854_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_855_ce = 1'b1;
    end else begin
        grp_fu_855_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_856_ce = 1'b1;
    end else begin
        grp_fu_856_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_857_ce = 1'b1;
    end else begin
        grp_fu_857_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_858_ce = 1'b1;
    end else begin
        grp_fu_858_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_859_ce = 1'b1;
    end else begin
        grp_fu_859_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_860_ce = 1'b1;
    end else begin
        grp_fu_860_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_861_ce = 1'b1;
    end else begin
        grp_fu_861_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_862_ce = 1'b1;
    end else begin
        grp_fu_862_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_863_ce = 1'b1;
    end else begin
        grp_fu_863_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_864_ce = 1'b1;
    end else begin
        grp_fu_864_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_866_ce = 1'b1;
    end else begin
        grp_fu_866_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_867_ce = 1'b1;
    end else begin
        grp_fu_867_ce = 1'b0;
    end
end

assign add_ln1118_1_fu_17671_p2 = ((sext_ln1118_76_fu_17661_p1) + (shl_ln1118_6_fu_17664_p3));

assign add_ln1118_2_fu_17735_p2 = ((shl_ln1118_7_fu_17717_p3) + (sext_ln1118_80_fu_17731_p1));

assign add_ln1118_fu_17625_p2 = ((shl_ln_fu_17607_p3) + (sext_ln1118_73_fu_17621_p1));

assign add_ln703_36_fu_17926_p2 = (trunc_ln708_31_reg_18953 + 16'd2428);

assign add_ln703_37_fu_17931_p2 = ((trunc_ln708_32_reg_18958) + (16'd63557));

assign add_ln703_38_fu_17936_p2 = (trunc_ln708_s_reg_18963 + 16'd2668);

assign add_ln703_39_fu_17941_p2 = (trunc_ln708_33_reg_18968 + 16'd770);

assign add_ln703_40_fu_17946_p2 = ((trunc_ln708_34_reg_18973) + (16'd65261));

assign add_ln703_41_fu_17951_p2 = (trunc_ln708_35_reg_18978 + 16'd1774);

assign add_ln703_42_fu_17956_p2 = ((trunc_ln708_36_reg_18983) + (16'd61620));

assign add_ln703_43_fu_17961_p2 = (trunc_ln708_37_reg_18988 + 16'd1134);

assign add_ln703_44_fu_17966_p2 = (trunc_ln708_38_reg_18993 + 16'd3344);

assign add_ln703_45_fu_17971_p2 = (trunc_ln708_39_reg_18998 + 16'd476);

assign add_ln703_46_fu_17976_p2 = ((trunc_ln708_40_reg_19003) + (16'd65055));

assign add_ln703_47_fu_17981_p2 = ((trunc_ln708_41_reg_19008) + (16'd63350));

assign add_ln703_48_fu_17986_p2 = (trunc_ln708_42_reg_19013 + 16'd6336);

assign add_ln703_49_fu_17991_p2 = (trunc_ln708_43_reg_19018 + 16'd779);

assign add_ln703_50_fu_17996_p2 = ((trunc_ln708_44_reg_19023) + (16'd65093));

assign add_ln703_51_fu_18001_p2 = ((trunc_ln708_45_reg_19028) + (16'd64452));

assign add_ln703_52_fu_18006_p2 = (trunc_ln708_46_reg_19033 + 16'd150);

assign add_ln703_53_fu_18011_p2 = ((trunc_ln708_47_reg_19038) + (16'd64356));

assign add_ln703_54_fu_18016_p2 = ((trunc_ln708_48_reg_19043) + (16'd61833));

assign add_ln703_55_fu_18021_p2 = ((trunc_ln708_49_reg_19048) + (16'd62693));

assign add_ln703_56_fu_18026_p2 = ((trunc_ln708_50_reg_19053) + (16'd65182));

assign add_ln703_57_fu_18031_p2 = ((trunc_ln708_51_reg_19058) + (16'd65467));

assign add_ln703_58_fu_18036_p2 = ((trunc_ln708_52_reg_19063) + (16'd65273));

assign add_ln703_59_fu_18041_p2 = ((trunc_ln708_53_reg_19068) + (16'd64093));

assign add_ln703_60_fu_18046_p2 = (trunc_ln708_54_reg_19073 + 16'd639);

assign add_ln703_61_fu_18051_p2 = ((trunc_ln708_55_reg_19078) + (16'd61811));

assign add_ln703_62_fu_18056_p2 = (trunc_ln708_56_reg_19083 + 16'd2997);

assign add_ln703_63_fu_18061_p2 = ((trunc_ln708_57_reg_19088) + (16'd65397));

assign add_ln703_64_fu_18066_p2 = ((trunc_ln708_58_reg_19093) + (16'd62604));

assign add_ln703_65_fu_18071_p2 = ((trunc_ln708_59_reg_19098) + (16'd60961));

assign add_ln703_66_fu_18076_p2 = (trunc_ln708_60_reg_19103 + 16'd3539);

assign add_ln703_67_fu_18081_p2 = ((trunc_ln708_61_reg_19108) + (16'd64305));

assign add_ln703_68_fu_18086_p2 = ((trunc_ln708_62_reg_19113) + (16'd64971));

assign add_ln703_69_fu_18091_p2 = (trunc_ln708_63_reg_19118 + 16'd427);

assign add_ln703_70_fu_18096_p2 = (trunc_ln708_64_reg_19123 + 16'd942);

assign add_ln703_71_fu_18101_p2 = ((trunc_ln708_65_reg_19128) + (16'd64448));

assign add_ln703_72_fu_18106_p2 = ((trunc_ln708_66_reg_19133) + (16'd61149));

assign add_ln703_73_fu_18111_p2 = ((trunc_ln708_67_reg_19138) + (16'd63555));

assign add_ln703_74_fu_18116_p2 = ((trunc_ln708_68_reg_19143) + (16'd64965));

assign add_ln703_75_fu_18121_p2 = ((trunc_ln708_69_reg_19148) + (16'd65184));

assign add_ln703_76_fu_18126_p2 = ((trunc_ln708_70_reg_19153) + (16'd65085));

assign add_ln703_77_fu_18131_p2 = ((trunc_ln708_71_reg_19158) + (16'd63019));

assign add_ln703_78_fu_18136_p2 = (trunc_ln708_72_reg_19163 + 16'd436);

assign add_ln703_79_fu_18141_p2 = ((trunc_ln708_73_reg_19168) + (16'd62012));

assign add_ln703_80_fu_18146_p2 = (trunc_ln708_74_reg_19173 + 16'd946);

assign add_ln703_81_fu_18151_p2 = ((trunc_ln708_75_reg_19178) + (16'd65281));

assign add_ln703_82_fu_18156_p2 = (trunc_ln708_76_reg_19183 + 16'd473);

assign add_ln703_83_fu_18161_p2 = ((trunc_ln708_77_reg_19188) + (16'd64458));

assign add_ln703_84_fu_18166_p2 = ((trunc_ln708_78_reg_19193) + (16'd65219));

assign add_ln703_85_fu_18171_p2 = (trunc_ln708_79_reg_19198 + 16'd1658);

assign add_ln703_86_fu_18176_p2 = (trunc_ln708_80_reg_19203 + 16'd2181);

assign add_ln703_87_fu_18181_p2 = (trunc_ln708_81_reg_19208 + 16'd1895);

assign add_ln703_88_fu_18186_p2 = (trunc_ln708_82_reg_19213 + 16'd792);

assign add_ln703_89_fu_18191_p2 = ((trunc_ln708_83_reg_19218) + (16'd62636));

assign add_ln703_90_fu_18196_p2 = (trunc_ln708_84_reg_19223 + 16'd1428);

assign add_ln703_91_fu_18201_p2 = ((trunc_ln708_85_reg_19228) + (16'd64938));

assign add_ln703_92_fu_18206_p2 = (trunc_ln708_86_reg_19233 + 16'd931);

assign add_ln703_93_fu_18211_p2 = ((trunc_ln708_87_reg_19238) + (16'd63398));

assign add_ln703_94_fu_18216_p2 = (trunc_ln708_88_reg_19243 + 16'd1118);

assign add_ln703_95_fu_18221_p2 = (trunc_ln708_89_reg_19248 + 16'd139);

assign add_ln703_96_fu_18226_p2 = (trunc_ln708_90_reg_19253 + 16'd1493);

assign add_ln703_97_fu_18231_p2 = (trunc_ln708_91_reg_19258 + 16'd396);

assign add_ln703_98_fu_18236_p2 = ((trunc_ln708_92_reg_19263) + (16'd61920));

assign add_ln703_fu_17921_p2 = ((trunc_ln_reg_18948) + (16'd64219));

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign grp_fu_804_p1 = 26'd1206;

assign grp_fu_805_p1 = 26'd1155;

assign grp_fu_806_p1 = 26'd1317;

assign grp_fu_807_p1 = 26'd1776;

assign grp_fu_808_p1 = 26'd753;

assign grp_fu_809_p1 = 26'd689;

assign grp_fu_810_p1 = 26'd1209;

assign grp_fu_811_p1 = 26'd880;

assign grp_fu_812_p1 = 26'd1483;

assign grp_fu_813_p1 = 26'd2953;

assign grp_fu_814_p1 = 26'd1379;

assign grp_fu_815_p1 = 26'd1208;

assign grp_fu_816_p1 = 26'd1089;

assign grp_fu_818_p1 = 26'd1827;

assign grp_fu_819_p1 = 26'd811;

assign grp_fu_820_p1 = 26'd1718;

assign grp_fu_821_p1 = 26'd1103;

assign grp_fu_822_p1 = 26'd1465;

assign grp_fu_823_p1 = 26'd1094;

assign grp_fu_824_p1 = 26'd1816;

assign grp_fu_825_p1 = 26'd850;

assign grp_fu_826_p1 = 26'd1241;

assign grp_fu_827_p1 = 26'd1315;

assign grp_fu_828_p1 = 26'd929;

assign grp_fu_829_p1 = 26'd931;

assign grp_fu_830_p1 = 26'd1361;

assign grp_fu_831_p1 = 26'd793;

assign grp_fu_832_p1 = 26'd999;

assign grp_fu_833_p1 = 26'd1589;

assign grp_fu_834_p1 = 26'd667;

assign grp_fu_835_p1 = 26'd1731;

assign grp_fu_837_p1 = 26'd1192;

assign grp_fu_838_p1 = 26'd2114;

assign grp_fu_839_p1 = 26'd832;

assign grp_fu_840_p1 = 26'd1254;

assign grp_fu_841_p1 = 26'd998;

assign grp_fu_842_p1 = 26'd1583;

assign grp_fu_843_p1 = 26'd947;

assign grp_fu_844_p1 = 26'd882;

assign grp_fu_845_p1 = 26'd936;

assign grp_fu_846_p1 = 26'd1168;

assign grp_fu_847_p1 = 26'd1604;

assign grp_fu_848_p1 = 26'd991;

assign grp_fu_849_p1 = 26'd1117;

assign grp_fu_850_p1 = 26'd817;

assign grp_fu_851_p1 = 26'd1116;

assign grp_fu_852_p1 = 26'd1611;

assign grp_fu_853_p1 = 26'd773;

assign grp_fu_854_p1 = 26'd2327;

assign grp_fu_855_p1 = 26'd1031;

assign grp_fu_856_p1 = 26'd868;

assign grp_fu_857_p1 = 26'd1751;

assign grp_fu_858_p1 = 26'd669;

assign grp_fu_859_p1 = 26'd1054;

assign grp_fu_860_p1 = 26'd1055;

assign grp_fu_861_p1 = 26'd1256;

assign grp_fu_862_p1 = 26'd1713;

assign grp_fu_863_p1 = 26'd1267;

assign grp_fu_864_p1 = 26'd901;

assign grp_fu_866_p1 = 26'd1881;

assign grp_fu_867_p1 = 26'd2145;

assign sext_ln1118_73_fu_17621_p1 = (shl_ln1118_5_fu_17614_p3);

assign sext_ln1118_76_fu_17661_p1 = data_42_V_read_2_reg_18631;

assign sext_ln1118_80_fu_17731_p1 = (shl_ln1118_8_fu_17724_p3);

assign shl_ln1118_5_fu_17614_p3 = {{data_39_V_read_2_reg_18637}, {7'd0}};

assign shl_ln1118_6_fu_17664_p3 = {{data_42_V_read_2_reg_18631}, {10'd0}};

assign shl_ln1118_7_fu_17717_p3 = {{data_46_V_read_2_reg_18625}, {10'd0}};

assign shl_ln1118_8_fu_17724_p3 = {{data_46_V_read_2_reg_18625}, {6'd0}};

assign shl_ln_fu_17607_p3 = {{data_39_V_read_2_reg_18637}, {10'd0}};

endmodule //normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;

wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [14:0] trunc_ln708_13_reg_5613;
reg   [14:0] trunc_ln708_13_reg_5613_pp0_iter1_reg;
reg   [13:0] tmp_385_reg_5703;
reg   [14:0] trunc_ln708_s_reg_5708;
reg   [15:0] trunc_ln708_4_reg_5713;
reg   [14:0] trunc_ln708_5_reg_5718;
reg   [15:0] trunc_ln708_6_reg_5723;
reg   [15:0] trunc_ln708_7_reg_5728;
reg   [14:0] trunc_ln708_8_reg_5733;
reg   [14:0] trunc_ln708_9_reg_5738;
reg   [15:0] trunc_ln708_1_reg_5743;
reg   [15:0] trunc_ln708_2_reg_5748;
reg   [15:0] trunc_ln708_3_reg_5753;
reg   [15:0] trunc_ln708_10_reg_5758;
reg   [15:0] trunc_ln708_11_reg_5763;
reg   [15:0] trunc_ln708_12_reg_5768;
reg   [15:0] trunc_ln708_14_reg_5773;
reg   [14:0] trunc_ln708_15_reg_5778;
reg   [14:0] trunc_ln708_16_reg_5783;
reg   [15:0] trunc_ln708_17_reg_5788;
reg   [14:0] trunc_ln708_18_reg_5793;
reg   [15:0] trunc_ln708_19_reg_5798;
reg   [15:0] trunc_ln708_20_reg_5803;
reg   [15:0] trunc_ln708_21_reg_5808;
reg   [15:0] trunc_ln708_22_reg_5813;
reg   [15:0] trunc_ln708_23_reg_5818;
reg   [15:0] trunc_ln708_24_reg_5823;
reg   [15:0] trunc_ln708_25_reg_5828;
reg   [15:0] trunc_ln708_26_reg_5833;
reg   [15:0] trunc_ln708_27_reg_5838;
reg   [15:0] trunc_ln708_28_reg_5843;
reg   [15:0] trunc_ln708_29_reg_5848;
reg   [14:0] trunc_ln708_30_reg_5853;
wire   [9:0] grp_fu_424_p1;
wire    ap_block_pp0_stage0;
wire   [9:0] grp_fu_425_p1;
wire   [8:0] grp_fu_426_p1;
wire   [8:0] grp_fu_427_p1;
wire   [9:0] grp_fu_428_p1;
wire   [9:0] grp_fu_429_p1;
wire   [8:0] grp_fu_430_p1;
wire   [9:0] grp_fu_431_p1;
wire   [8:0] grp_fu_432_p1;
wire   [8:0] grp_fu_433_p1;
wire   [9:0] grp_fu_435_p1;
wire   [7:0] grp_fu_436_p1;
wire   [9:0] grp_fu_437_p1;
wire   [8:0] grp_fu_438_p1;
wire   [8:0] grp_fu_439_p1;
wire   [9:0] grp_fu_440_p1;
wire   [9:0] grp_fu_441_p1;
wire   [9:0] grp_fu_442_p1;
wire   [9:0] grp_fu_443_p1;
wire   [10:0] grp_fu_444_p1;
wire   [8:0] grp_fu_445_p1;
wire   [10:0] grp_fu_446_p1;
wire   [9:0] grp_fu_447_p1;
wire   [9:0] grp_fu_448_p1;
wire   [10:0] grp_fu_449_p1;
wire   [9:0] grp_fu_450_p1;
wire   [9:0] grp_fu_451_p1;
wire   [9:0] grp_fu_452_p1;
wire   [9:0] grp_fu_453_p1;
wire   [9:0] grp_fu_454_p1;
wire   [9:0] grp_fu_455_p1;
wire   [23:0] shl_ln_fu_4712_p3;
wire   [16:0] shl_ln1118_9_fu_4724_p3;
wire   [24:0] sext_ln1118_17_fu_4720_p1;
wire   [24:0] sext_ln1118_18_fu_4732_p1;
wire   [24:0] sub_ln1118_fu_4736_p2;
wire   [23:0] grp_fu_436_p2;
wire   [24:0] grp_fu_426_p2;
wire   [25:0] grp_fu_435_p2;
wire   [24:0] grp_fu_439_p2;
wire   [25:0] grp_fu_440_p2;
wire   [25:0] grp_fu_449_p2;
wire   [24:0] grp_fu_432_p2;
wire   [24:0] grp_fu_430_p2;
wire   [25:0] grp_fu_441_p2;
wire   [25:0] grp_fu_451_p2;
wire   [25:0] grp_fu_425_p2;
wire   [25:0] grp_fu_450_p2;
wire   [25:0] grp_fu_428_p2;
wire   [25:0] grp_fu_442_p2;
wire   [25:0] grp_fu_446_p2;
wire   [24:0] grp_fu_427_p2;
wire   [24:0] grp_fu_445_p2;
wire   [25:0] grp_fu_424_p2;
wire   [24:0] grp_fu_438_p2;
wire   [25:0] grp_fu_453_p2;
wire   [25:0] grp_fu_431_p2;
wire   [25:0] grp_fu_429_p2;
wire   [25:0] grp_fu_455_p2;
wire   [25:0] grp_fu_444_p2;
wire   [25:0] grp_fu_448_p2;
wire   [25:0] grp_fu_443_p2;
wire   [25:0] grp_fu_452_p2;
wire   [25:0] grp_fu_437_p2;
wire   [25:0] grp_fu_447_p2;
wire   [25:0] grp_fu_454_p2;
wire   [24:0] grp_fu_433_p2;
wire   [14:0] sext_ln703_fu_5147_p1;
wire   [14:0] add_ln703_fu_5150_p2;
wire   [15:0] sext_ln708_fu_5160_p1;
wire   [15:0] sext_ln708_4_fu_5174_p1;
wire   [15:0] sext_ln708_5_fu_5193_p1;
wire   [15:0] sext_ln708_6_fu_5202_p1;
wire   [15:0] sext_ln708_7_fu_5241_p1;
wire   [15:0] sext_ln708_8_fu_5255_p1;
wire   [15:0] sext_ln708_9_fu_5264_p1;
wire   [15:0] sext_ln708_10_fu_5278_p1;
wire   [15:0] sext_ln708_11_fu_5342_p1;
wire   [15:0] sext_ln703_2_fu_5156_p1;
wire   [15:0] add_ln703_5_fu_5163_p2;
wire   [15:0] add_ln703_6_fu_5169_p2;
wire   [15:0] add_ln703_7_fu_5177_p2;
wire   [15:0] add_ln703_8_fu_5183_p2;
wire   [15:0] add_ln703_9_fu_5188_p2;
wire   [15:0] add_ln703_10_fu_5196_p2;
wire   [15:0] add_ln703_11_fu_5205_p2;
wire   [15:0] add_ln703_12_fu_5211_p2;
wire   [15:0] add_ln703_13_fu_5216_p2;
wire   [15:0] add_ln703_14_fu_5221_p2;
wire   [15:0] add_ln703_15_fu_5226_p2;
wire   [15:0] add_ln703_16_fu_5231_p2;
wire   [15:0] add_ln703_17_fu_5236_p2;
wire   [15:0] add_ln703_18_fu_5244_p2;
wire   [15:0] add_ln703_19_fu_5250_p2;
wire   [15:0] add_ln703_20_fu_5258_p2;
wire   [15:0] add_ln703_21_fu_5267_p2;
wire   [15:0] add_ln703_22_fu_5273_p2;
wire   [15:0] add_ln703_23_fu_5281_p2;
wire   [15:0] add_ln703_24_fu_5287_p2;
wire   [15:0] add_ln703_25_fu_5292_p2;
wire   [15:0] add_ln703_26_fu_5297_p2;
wire   [15:0] add_ln703_27_fu_5302_p2;
wire   [15:0] add_ln703_28_fu_5307_p2;
wire   [15:0] add_ln703_29_fu_5312_p2;
wire   [15:0] add_ln703_30_fu_5317_p2;
wire   [15:0] add_ln703_31_fu_5322_p2;
wire   [15:0] add_ln703_32_fu_5327_p2;
wire   [15:0] add_ln703_33_fu_5332_p2;
wire   [15:0] add_ln703_34_fu_5337_p2;
wire   [15:0] add_ln703_35_fu_5345_p2;
reg    grp_fu_424_ce;
reg    grp_fu_425_ce;
reg    grp_fu_426_ce;
reg    grp_fu_427_ce;
reg    grp_fu_428_ce;
reg    grp_fu_429_ce;
reg    grp_fu_430_ce;
reg    grp_fu_431_ce;
reg    grp_fu_432_ce;
reg    grp_fu_433_ce;
reg    grp_fu_435_ce;
reg    grp_fu_436_ce;
reg    grp_fu_437_ce;
reg    grp_fu_438_ce;
reg    grp_fu_439_ce;
reg    grp_fu_440_ce;
reg    grp_fu_441_ce;
reg    grp_fu_442_ce;
reg    grp_fu_443_ce;
reg    grp_fu_444_ce;
reg    grp_fu_445_ce;
reg    grp_fu_446_ce;
reg    grp_fu_447_ce;
reg    grp_fu_448_ce;
reg    grp_fu_449_ce;
reg    grp_fu_450_ce;
reg    grp_fu_451_ce;
reg    grp_fu_452_ce;
reg    grp_fu_453_ce;
reg    grp_fu_454_ce;
reg    grp_fu_455_ce;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U385(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_18_V_read_int_reg),
    .din1(grp_fu_424_p1),
    .ce(grp_fu_424_ce),
    .dout(grp_fu_424_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U386(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_10_V_read_int_reg),
    .din1(grp_fu_425_p1),
    .ce(grp_fu_425_ce),
    .dout(grp_fu_425_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U387(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_1_V_read_int_reg),
    .din1(grp_fu_426_p1),
    .ce(grp_fu_426_ce),
    .dout(grp_fu_426_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U388(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_16_V_read_int_reg),
    .din1(grp_fu_427_p1),
    .ce(grp_fu_427_ce),
    .dout(grp_fu_427_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U389(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_12_V_read_int_reg),
    .din1(grp_fu_428_p1),
    .ce(grp_fu_428_ce),
    .dout(grp_fu_428_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U390(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_22_V_read_int_reg),
    .din1(grp_fu_429_p1),
    .ce(grp_fu_429_ce),
    .dout(grp_fu_429_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U391(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_7_V_read_int_reg),
    .din1(grp_fu_430_p1),
    .ce(grp_fu_430_ce),
    .dout(grp_fu_430_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U392(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_21_V_read_int_reg),
    .din1(grp_fu_431_p1),
    .ce(grp_fu_431_ce),
    .dout(grp_fu_431_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U393(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_6_V_read_int_reg),
    .din1(grp_fu_432_p1),
    .ce(grp_fu_432_ce),
    .dout(grp_fu_432_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U394(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_31_V_read_int_reg),
    .din1(grp_fu_433_p1),
    .ce(grp_fu_433_ce),
    .dout(grp_fu_433_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U395(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_2_V_read_int_reg),
    .din1(grp_fu_435_p1),
    .ce(grp_fu_435_ce),
    .dout(grp_fu_435_p2)
);

myproject_mul_16s_8ns_24_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 24 ))
myproject_mul_16s_8ns_24_2_0_U396(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_0_V_read_int_reg),
    .din1(grp_fu_436_p1),
    .ce(grp_fu_436_ce),
    .dout(grp_fu_436_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U397(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_28_V_read_int_reg),
    .din1(grp_fu_437_p1),
    .ce(grp_fu_437_ce),
    .dout(grp_fu_437_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U398(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_19_V_read_int_reg),
    .din1(grp_fu_438_p1),
    .ce(grp_fu_438_ce),
    .dout(grp_fu_438_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U399(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_3_V_read_int_reg),
    .din1(grp_fu_439_p1),
    .ce(grp_fu_439_ce),
    .dout(grp_fu_439_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U400(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_4_V_read_int_reg),
    .din1(grp_fu_440_p1),
    .ce(grp_fu_440_ce),
    .dout(grp_fu_440_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U401(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_8_V_read_int_reg),
    .din1(grp_fu_441_p1),
    .ce(grp_fu_441_ce),
    .dout(grp_fu_441_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U402(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_13_V_read_int_reg),
    .din1(grp_fu_442_p1),
    .ce(grp_fu_442_ce),
    .dout(grp_fu_442_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U403(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_26_V_read_int_reg),
    .din1(grp_fu_443_p1),
    .ce(grp_fu_443_ce),
    .dout(grp_fu_443_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U404(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_24_V_read_int_reg),
    .din1(grp_fu_444_p1),
    .ce(grp_fu_444_ce),
    .dout(grp_fu_444_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U405(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_17_V_read_int_reg),
    .din1(grp_fu_445_p1),
    .ce(grp_fu_445_ce),
    .dout(grp_fu_445_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U406(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_15_V_read_int_reg),
    .din1(grp_fu_446_p1),
    .ce(grp_fu_446_ce),
    .dout(grp_fu_446_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U407(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_29_V_read_int_reg),
    .din1(grp_fu_447_p1),
    .ce(grp_fu_447_ce),
    .dout(grp_fu_447_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U408(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_25_V_read_int_reg),
    .din1(grp_fu_448_p1),
    .ce(grp_fu_448_ce),
    .dout(grp_fu_448_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U409(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_5_V_read_int_reg),
    .din1(grp_fu_449_p1),
    .ce(grp_fu_449_ce),
    .dout(grp_fu_449_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U410(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_11_V_read_int_reg),
    .din1(grp_fu_450_p1),
    .ce(grp_fu_450_ce),
    .dout(grp_fu_450_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U411(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_9_V_read_int_reg),
    .din1(grp_fu_451_p1),
    .ce(grp_fu_451_ce),
    .dout(grp_fu_451_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U412(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_27_V_read_int_reg),
    .din1(grp_fu_452_p1),
    .ce(grp_fu_452_ce),
    .dout(grp_fu_452_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U413(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_20_V_read_int_reg),
    .din1(grp_fu_453_p1),
    .ce(grp_fu_453_ce),
    .dout(grp_fu_453_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U414(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_30_V_read_int_reg),
    .din1(grp_fu_454_p1),
    .ce(grp_fu_454_ce),
    .dout(grp_fu_454_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U415(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_23_V_read_int_reg),
    .din1(grp_fu_455_p1),
    .ce(grp_fu_455_ce),
    .dout(grp_fu_455_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= sext_ln703_2_fu_5156_p1;
        ap_return_10_int_reg <= add_ln703_14_fu_5221_p2;
        ap_return_11_int_reg <= add_ln703_15_fu_5226_p2;
        ap_return_12_int_reg <= add_ln703_16_fu_5231_p2;
        ap_return_13_int_reg <= add_ln703_17_fu_5236_p2;
        ap_return_14_int_reg <= add_ln703_18_fu_5244_p2;
        ap_return_15_int_reg <= add_ln703_19_fu_5250_p2;
        ap_return_16_int_reg <= add_ln703_20_fu_5258_p2;
        ap_return_17_int_reg <= add_ln703_21_fu_5267_p2;
        ap_return_18_int_reg <= add_ln703_22_fu_5273_p2;
        ap_return_19_int_reg <= add_ln703_23_fu_5281_p2;
        ap_return_1_int_reg <= add_ln703_5_fu_5163_p2;
        ap_return_20_int_reg <= add_ln703_24_fu_5287_p2;
        ap_return_21_int_reg <= add_ln703_25_fu_5292_p2;
        ap_return_22_int_reg <= add_ln703_26_fu_5297_p2;
        ap_return_23_int_reg <= add_ln703_27_fu_5302_p2;
        ap_return_24_int_reg <= add_ln703_28_fu_5307_p2;
        ap_return_25_int_reg <= add_ln703_29_fu_5312_p2;
        ap_return_26_int_reg <= add_ln703_30_fu_5317_p2;
        ap_return_27_int_reg <= add_ln703_31_fu_5322_p2;
        ap_return_28_int_reg <= add_ln703_32_fu_5327_p2;
        ap_return_29_int_reg <= add_ln703_33_fu_5332_p2;
        ap_return_2_int_reg <= add_ln703_6_fu_5169_p2;
        ap_return_30_int_reg <= add_ln703_34_fu_5337_p2;
        ap_return_31_int_reg <= add_ln703_35_fu_5345_p2;
        ap_return_3_int_reg <= add_ln703_7_fu_5177_p2;
        ap_return_4_int_reg <= add_ln703_8_fu_5183_p2;
        ap_return_5_int_reg <= add_ln703_9_fu_5188_p2;
        ap_return_6_int_reg <= add_ln703_10_fu_5196_p2;
        ap_return_7_int_reg <= add_ln703_11_fu_5205_p2;
        ap_return_8_int_reg <= add_ln703_12_fu_5211_p2;
        ap_return_9_int_reg <= add_ln703_13_fu_5216_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        tmp_385_reg_5703 <= {{grp_fu_436_p2[23:10]}};
        trunc_ln708_10_reg_5758 <= {{grp_fu_450_p2[25:10]}};
        trunc_ln708_11_reg_5763 <= {{grp_fu_428_p2[25:10]}};
        trunc_ln708_12_reg_5768 <= {{grp_fu_442_p2[25:10]}};
        trunc_ln708_13_reg_5613 <= {{sub_ln1118_fu_4736_p2[24:10]}};
        trunc_ln708_13_reg_5613_pp0_iter1_reg <= trunc_ln708_13_reg_5613;
        trunc_ln708_14_reg_5773 <= {{grp_fu_446_p2[25:10]}};
        trunc_ln708_15_reg_5778 <= {{grp_fu_427_p2[24:10]}};
        trunc_ln708_16_reg_5783 <= {{grp_fu_445_p2[24:10]}};
        trunc_ln708_17_reg_5788 <= {{grp_fu_424_p2[25:10]}};
        trunc_ln708_18_reg_5793 <= {{grp_fu_438_p2[24:10]}};
        trunc_ln708_19_reg_5798 <= {{grp_fu_453_p2[25:10]}};
        trunc_ln708_1_reg_5743 <= {{grp_fu_441_p2[25:10]}};
        trunc_ln708_20_reg_5803 <= {{grp_fu_431_p2[25:10]}};
        trunc_ln708_21_reg_5808 <= {{grp_fu_429_p2[25:10]}};
        trunc_ln708_22_reg_5813 <= {{grp_fu_455_p2[25:10]}};
        trunc_ln708_23_reg_5818 <= {{grp_fu_444_p2[25:10]}};
        trunc_ln708_24_reg_5823 <= {{grp_fu_448_p2[25:10]}};
        trunc_ln708_25_reg_5828 <= {{grp_fu_443_p2[25:10]}};
        trunc_ln708_26_reg_5833 <= {{grp_fu_452_p2[25:10]}};
        trunc_ln708_27_reg_5838 <= {{grp_fu_437_p2[25:10]}};
        trunc_ln708_28_reg_5843 <= {{grp_fu_447_p2[25:10]}};
        trunc_ln708_29_reg_5848 <= {{grp_fu_454_p2[25:10]}};
        trunc_ln708_2_reg_5748 <= {{grp_fu_451_p2[25:10]}};
        trunc_ln708_30_reg_5853 <= {{grp_fu_433_p2[24:10]}};
        trunc_ln708_3_reg_5753 <= {{grp_fu_425_p2[25:10]}};
        trunc_ln708_4_reg_5713 <= {{grp_fu_435_p2[25:10]}};
        trunc_ln708_5_reg_5718 <= {{grp_fu_439_p2[24:10]}};
        trunc_ln708_6_reg_5723 <= {{grp_fu_440_p2[25:10]}};
        trunc_ln708_7_reg_5728 <= {{grp_fu_449_p2[25:10]}};
        trunc_ln708_8_reg_5733 <= {{grp_fu_432_p2[24:10]}};
        trunc_ln708_9_reg_5738 <= {{grp_fu_430_p2[24:10]}};
        trunc_ln708_s_reg_5708 <= {{grp_fu_426_p2[24:10]}};
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = sext_ln703_2_fu_5156_p1;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = add_ln703_5_fu_5163_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = add_ln703_14_fu_5221_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = add_ln703_15_fu_5226_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = add_ln703_16_fu_5231_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = add_ln703_17_fu_5236_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = add_ln703_18_fu_5244_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = add_ln703_19_fu_5250_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = add_ln703_20_fu_5258_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = add_ln703_21_fu_5267_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = add_ln703_22_fu_5273_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = add_ln703_23_fu_5281_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = add_ln703_6_fu_5169_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = add_ln703_24_fu_5287_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = add_ln703_25_fu_5292_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = add_ln703_26_fu_5297_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = add_ln703_27_fu_5302_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = add_ln703_28_fu_5307_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = add_ln703_29_fu_5312_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = add_ln703_30_fu_5317_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = add_ln703_31_fu_5322_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = add_ln703_32_fu_5327_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = add_ln703_33_fu_5332_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = add_ln703_7_fu_5177_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = add_ln703_34_fu_5337_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = add_ln703_35_fu_5345_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = add_ln703_8_fu_5183_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = add_ln703_9_fu_5188_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = add_ln703_10_fu_5196_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = add_ln703_11_fu_5205_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = add_ln703_12_fu_5211_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = add_ln703_13_fu_5216_p2;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_424_ce = 1'b1;
    end else begin
        grp_fu_424_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_425_ce = 1'b1;
    end else begin
        grp_fu_425_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_426_ce = 1'b1;
    end else begin
        grp_fu_426_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_427_ce = 1'b1;
    end else begin
        grp_fu_427_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_428_ce = 1'b1;
    end else begin
        grp_fu_428_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_429_ce = 1'b1;
    end else begin
        grp_fu_429_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_430_ce = 1'b1;
    end else begin
        grp_fu_430_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_431_ce = 1'b1;
    end else begin
        grp_fu_431_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_432_ce = 1'b1;
    end else begin
        grp_fu_432_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_433_ce = 1'b1;
    end else begin
        grp_fu_433_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_435_ce = 1'b1;
    end else begin
        grp_fu_435_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_436_ce = 1'b1;
    end else begin
        grp_fu_436_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_437_ce = 1'b1;
    end else begin
        grp_fu_437_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_438_ce = 1'b1;
    end else begin
        grp_fu_438_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_439_ce = 1'b1;
    end else begin
        grp_fu_439_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_440_ce = 1'b1;
    end else begin
        grp_fu_440_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_441_ce = 1'b1;
    end else begin
        grp_fu_441_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_442_ce = 1'b1;
    end else begin
        grp_fu_442_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_443_ce = 1'b1;
    end else begin
        grp_fu_443_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_444_ce = 1'b1;
    end else begin
        grp_fu_444_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_445_ce = 1'b1;
    end else begin
        grp_fu_445_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_446_ce = 1'b1;
    end else begin
        grp_fu_446_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_447_ce = 1'b1;
    end else begin
        grp_fu_447_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_448_ce = 1'b1;
    end else begin
        grp_fu_448_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_449_ce = 1'b1;
    end else begin
        grp_fu_449_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_450_ce = 1'b1;
    end else begin
        grp_fu_450_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_451_ce = 1'b1;
    end else begin
        grp_fu_451_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_452_ce = 1'b1;
    end else begin
        grp_fu_452_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_453_ce = 1'b1;
    end else begin
        grp_fu_453_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_454_ce = 1'b1;
    end else begin
        grp_fu_454_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_455_ce = 1'b1;
    end else begin
        grp_fu_455_ce = 1'b0;
    end
end

assign add_ln703_10_fu_5196_p2 = ((sext_ln708_5_fu_5193_p1) + (16'd446));

assign add_ln703_11_fu_5205_p2 = ((sext_ln708_6_fu_5202_p1) + (16'd597));

assign add_ln703_12_fu_5211_p2 = (trunc_ln708_1_reg_5743 + 16'd408);

assign add_ln703_13_fu_5216_p2 = (trunc_ln708_2_reg_5748 + 16'd634);

assign add_ln703_14_fu_5221_p2 = ((trunc_ln708_3_reg_5753) + (16'd65224));

assign add_ln703_15_fu_5226_p2 = (trunc_ln708_10_reg_5758 + 16'd1821);

assign add_ln703_16_fu_5231_p2 = ((trunc_ln708_11_reg_5763) + (16'd64651));

assign add_ln703_17_fu_5236_p2 = (trunc_ln708_12_reg_5768 + 16'd672);

assign add_ln703_18_fu_5244_p2 = ((sext_ln708_7_fu_5241_p1) + (16'd445));

assign add_ln703_19_fu_5250_p2 = (trunc_ln708_14_reg_5773 + 16'd15);

assign add_ln703_20_fu_5258_p2 = ((sext_ln708_8_fu_5255_p1) + (16'd64909));

assign add_ln703_21_fu_5267_p2 = ((sext_ln708_9_fu_5264_p1) + (16'd65100));

assign add_ln703_22_fu_5273_p2 = ((trunc_ln708_17_reg_5788) + (16'd64899));

assign add_ln703_23_fu_5281_p2 = ((sext_ln708_10_fu_5278_p1) + (16'd439));

assign add_ln703_24_fu_5287_p2 = ((trunc_ln708_19_reg_5798) + (16'd64895));

assign add_ln703_25_fu_5292_p2 = (trunc_ln708_20_reg_5803 + 16'd379);

assign add_ln703_26_fu_5297_p2 = ((trunc_ln708_21_reg_5808) + (16'd65532));

assign add_ln703_27_fu_5302_p2 = ((trunc_ln708_22_reg_5813) + (16'd65400));

assign add_ln703_28_fu_5307_p2 = (trunc_ln708_23_reg_5818 + 16'd622);

assign add_ln703_29_fu_5312_p2 = (trunc_ln708_24_reg_5823 + 16'd15);

assign add_ln703_30_fu_5317_p2 = ((trunc_ln708_25_reg_5828) + (16'd65459));

assign add_ln703_31_fu_5322_p2 = (trunc_ln708_26_reg_5833 + 16'd416);

assign add_ln703_32_fu_5327_p2 = (trunc_ln708_27_reg_5838 + 16'd31);

assign add_ln703_33_fu_5332_p2 = ((trunc_ln708_28_reg_5843) + (16'd65502));

assign add_ln703_34_fu_5337_p2 = ((trunc_ln708_29_reg_5848) + (16'd64870));

assign add_ln703_35_fu_5345_p2 = ((sext_ln708_11_fu_5342_p1) + (16'd288));

assign add_ln703_5_fu_5163_p2 = ((sext_ln708_fu_5160_p1) + (16'd65252));

assign add_ln703_6_fu_5169_p2 = (trunc_ln708_4_reg_5713 + 16'd617);

assign add_ln703_7_fu_5177_p2 = ((sext_ln708_4_fu_5174_p1) + (16'd129));

assign add_ln703_8_fu_5183_p2 = ((trunc_ln708_6_reg_5723) + (16'd64666));

assign add_ln703_9_fu_5188_p2 = ((trunc_ln708_7_reg_5728) + (16'd65475));

assign add_ln703_fu_5150_p2 = ((sext_ln703_fu_5147_p1) + (15'd32383));

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign grp_fu_424_p1 = 26'd421;

assign grp_fu_425_p1 = 26'd353;

assign grp_fu_426_p1 = 25'd197;

assign grp_fu_427_p1 = 25'd198;

assign grp_fu_428_p1 = 26'd365;

assign grp_fu_429_p1 = 26'd359;

assign grp_fu_430_p1 = 25'd194;

assign grp_fu_431_p1 = 26'd358;

assign grp_fu_432_p1 = 25'd198;

assign grp_fu_433_p1 = 25'd253;

assign grp_fu_435_p1 = 26'd316;

assign grp_fu_436_p1 = 24'd125;

assign grp_fu_437_p1 = 26'd453;

assign grp_fu_438_p1 = 25'd233;

assign grp_fu_439_p1 = 25'd220;

assign grp_fu_440_p1 = 26'd341;

assign grp_fu_441_p1 = 26'd294;

assign grp_fu_442_p1 = 26'd310;

assign grp_fu_443_p1 = 26'd280;

assign grp_fu_444_p1 = 26'd617;

assign grp_fu_445_p1 = 25'd241;

assign grp_fu_446_p1 = 26'd618;

assign grp_fu_447_p1 = 26'd319;

assign grp_fu_448_p1 = 26'd385;

assign grp_fu_449_p1 = 26'd616;

assign grp_fu_450_p1 = 26'd486;

assign grp_fu_451_p1 = 26'd447;

assign grp_fu_452_p1 = 26'd324;

assign grp_fu_453_p1 = 26'd484;

assign grp_fu_454_p1 = 26'd487;

assign grp_fu_455_p1 = 26'd485;

assign sext_ln1118_17_fu_4720_p1 = (shl_ln_fu_4712_p3);

assign sext_ln1118_18_fu_4732_p1 = (shl_ln1118_9_fu_4724_p3);

assign sext_ln703_2_fu_5156_p1 = (add_ln703_fu_5150_p2);

assign sext_ln703_fu_5147_p1 = (tmp_385_reg_5703);

assign sext_ln708_10_fu_5278_p1 = (trunc_ln708_18_reg_5793);

assign sext_ln708_11_fu_5342_p1 = (trunc_ln708_30_reg_5853);

assign sext_ln708_4_fu_5174_p1 = (trunc_ln708_5_reg_5718);

assign sext_ln708_5_fu_5193_p1 = (trunc_ln708_8_reg_5733);

assign sext_ln708_6_fu_5202_p1 = (trunc_ln708_9_reg_5738);

assign sext_ln708_7_fu_5241_p1 = (trunc_ln708_13_reg_5613_pp0_iter1_reg);

assign sext_ln708_8_fu_5255_p1 = (trunc_ln708_15_reg_5778);

assign sext_ln708_9_fu_5264_p1 = (trunc_ln708_16_reg_5783);

assign sext_ln708_fu_5160_p1 = (trunc_ln708_s_reg_5708);

assign shl_ln1118_9_fu_4724_p3 = {{data_14_V_read_int_reg}, {1'd0}};

assign shl_ln_fu_4712_p3 = {{data_14_V_read_int_reg}, {8'd0}};

assign sub_ln1118_fu_4736_p2 = ((sext_ln1118_17_fu_4720_p1) - (sext_ln1118_18_fu_4732_p1));

endmodule //normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;

wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [14:0] trunc_ln708_22_reg_5489;
reg   [14:0] trunc_ln708_22_reg_5489_pp0_iter1_reg;
reg   [14:0] trunc_ln708_27_reg_5514;
reg   [14:0] trunc_ln708_27_reg_5514_pp0_iter1_reg;
reg   [13:0] tmp_386_reg_5519;
reg   [13:0] tmp_386_reg_5519_pp0_iter1_reg;
reg   [14:0] trunc_ln_reg_5539;
reg   [14:0] trunc_ln708_1_reg_5544;
reg   [14:0] trunc_ln708_2_reg_5549;
reg   [14:0] trunc_ln708_3_reg_5554;
reg   [14:0] trunc_ln708_4_reg_5559;
reg   [14:0] trunc_ln708_5_reg_5564;
reg   [15:0] trunc_ln708_6_reg_5569;
reg   [14:0] trunc_ln708_7_reg_5574;
reg   [14:0] trunc_ln708_8_reg_5579;
reg   [15:0] trunc_ln708_9_reg_5584;
reg   [14:0] trunc_ln708_10_reg_5589;
reg   [15:0] trunc_ln708_11_reg_5594;
reg   [14:0] trunc_ln708_12_reg_5599;
reg   [14:0] trunc_ln708_13_reg_5604;
reg   [14:0] trunc_ln708_14_reg_5609;
reg   [14:0] trunc_ln708_15_reg_5614;
reg   [15:0] trunc_ln708_16_reg_5619;
reg   [15:0] trunc_ln708_17_reg_5624;
reg   [14:0] trunc_ln708_18_reg_5629;
reg   [15:0] trunc_ln708_19_reg_5634;
reg   [14:0] trunc_ln708_20_reg_5639;
reg   [14:0] trunc_ln708_21_reg_5644;
reg   [14:0] trunc_ln708_23_reg_5649;
reg   [14:0] trunc_ln708_24_reg_5654;
reg   [14:0] trunc_ln708_25_reg_5659;
reg   [14:0] trunc_ln708_26_reg_5664;
reg   [14:0] trunc_ln708_29_reg_5669;
reg   [14:0] trunc_ln708_30_reg_5674;
reg   [15:0] trunc_ln708_31_reg_5679;
wire   [8:0] grp_fu_428_p1;
wire    ap_block_pp0_stage0;
wire   [8:0] grp_fu_430_p1;
wire   [8:0] grp_fu_431_p1;
wire   [8:0] grp_fu_432_p1;
wire   [8:0] grp_fu_433_p1;
wire   [8:0] grp_fu_435_p1;
wire   [8:0] grp_fu_436_p1;
wire   [9:0] grp_fu_437_p1;
wire   [9:0] grp_fu_438_p1;
wire   [9:0] grp_fu_439_p1;
wire   [9:0] grp_fu_440_p1;
wire   [8:0] grp_fu_441_p1;
wire   [8:0] grp_fu_442_p1;
wire   [8:0] grp_fu_443_p1;
wire   [8:0] grp_fu_444_p1;
wire   [9:0] grp_fu_445_p1;
wire   [8:0] grp_fu_446_p1;
wire   [8:0] grp_fu_447_p1;
wire   [8:0] grp_fu_448_p1;
wire   [8:0] grp_fu_449_p1;
wire   [8:0] grp_fu_451_p1;
wire   [8:0] grp_fu_452_p1;
wire   [9:0] grp_fu_453_p1;
wire   [8:0] grp_fu_454_p1;
wire   [9:0] grp_fu_455_p1;
wire   [8:0] grp_fu_456_p1;
wire   [8:0] grp_fu_457_p1;
wire   [8:0] grp_fu_458_p1;
wire   [8:0] grp_fu_459_p1;
wire   [15:0] sext_ln1118_22_fu_4486_p0;
wire   [15:0] shl_ln_fu_4490_p1;
wire   [23:0] shl_ln_fu_4490_p3;
wire   [24:0] sext_ln1118_23_fu_4498_p1;
wire   [24:0] sext_ln1118_22_fu_4486_p1;
wire   [24:0] add_ln1118_fu_4502_p2;
wire   [23:0] shl_ln1118_1_fu_4538_p3;
wire   [21:0] shl_ln1118_2_fu_4550_p3;
wire   [24:0] sext_ln1118_29_fu_4558_p1;
wire   [24:0] sext_ln1118_28_fu_4546_p1;
wire   [24:0] add_ln1118_1_fu_4562_p2;
wire   [22:0] shl_ln1118_3_fu_4578_p3;
wire   [20:0] shl_ln1118_4_fu_4590_p3;
wire   [23:0] sext_ln1118_31_fu_4598_p1;
wire   [23:0] sext_ln1118_30_fu_4586_p1;
wire   [23:0] add_ln1118_2_fu_4602_p2;
wire   [24:0] grp_fu_435_p2;
wire   [24:0] grp_fu_442_p2;
wire   [24:0] grp_fu_446_p2;
wire   [24:0] grp_fu_458_p2;
wire   [24:0] grp_fu_444_p2;
wire   [24:0] grp_fu_454_p2;
wire   [25:0] grp_fu_437_p2;
wire   [24:0] grp_fu_452_p2;
wire   [24:0] grp_fu_436_p2;
wire   [25:0] grp_fu_445_p2;
wire   [24:0] grp_fu_448_p2;
wire   [25:0] grp_fu_438_p2;
wire   [24:0] grp_fu_443_p2;
wire   [24:0] grp_fu_431_p2;
wire   [24:0] grp_fu_428_p2;
wire   [24:0] grp_fu_456_p2;
wire   [25:0] grp_fu_455_p2;
wire   [25:0] grp_fu_439_p2;
wire   [24:0] grp_fu_433_p2;
wire   [25:0] grp_fu_453_p2;
wire   [24:0] grp_fu_451_p2;
wire   [24:0] grp_fu_430_p2;
wire   [24:0] grp_fu_447_p2;
wire   [24:0] grp_fu_449_p2;
wire   [24:0] grp_fu_441_p2;
wire   [24:0] grp_fu_459_p2;
wire   [24:0] grp_fu_457_p2;
wire   [24:0] grp_fu_432_p2;
wire   [25:0] grp_fu_440_p2;
wire   [15:0] sext_ln708_fu_4923_p1;
wire   [15:0] sext_ln708_1_fu_4932_p1;
wire   [15:0] sext_ln708_2_fu_4941_p1;
wire   [15:0] sext_ln708_3_fu_4950_p1;
wire   [15:0] sext_ln708_4_fu_4959_p1;
wire   [15:0] sext_ln708_5_fu_4968_p1;
wire   [15:0] sext_ln708_6_fu_4982_p1;
wire   [15:0] sext_ln708_7_fu_4991_p1;
wire   [15:0] sext_ln708_8_fu_5005_p1;
wire   [15:0] sext_ln708_9_fu_5019_p1;
wire   [15:0] sext_ln708_10_fu_5028_p1;
wire   [15:0] sext_ln708_11_fu_5037_p1;
wire   [15:0] sext_ln708_12_fu_5046_p1;
wire   [15:0] sext_ln708_13_fu_5065_p1;
wire   [15:0] sext_ln708_14_fu_5079_p1;
wire   [15:0] sext_ln708_15_fu_5088_p1;
wire   [15:0] sext_ln708_16_fu_5097_p1;
wire   [15:0] sext_ln708_17_fu_5106_p1;
wire   [15:0] sext_ln708_18_fu_5115_p1;
wire   [15:0] sext_ln708_19_fu_5124_p1;
wire   [15:0] sext_ln708_20_fu_5133_p1;
wire   [15:0] sext_ln708_21_fu_5142_p1;
wire   [14:0] sext_ln703_fu_5151_p1;
wire   [14:0] add_ln703_126_fu_5154_p2;
wire   [15:0] sext_ln708_22_fu_5164_p1;
wire   [15:0] sext_ln708_23_fu_5173_p1;
wire   [15:0] add_ln703_fu_4926_p2;
wire   [15:0] add_ln703_99_fu_4935_p2;
wire   [15:0] add_ln703_100_fu_4944_p2;
wire   [15:0] add_ln703_101_fu_4953_p2;
wire   [15:0] add_ln703_102_fu_4962_p2;
wire   [15:0] add_ln703_103_fu_4971_p2;
wire   [15:0] add_ln703_104_fu_4977_p2;
wire   [15:0] add_ln703_105_fu_4985_p2;
wire   [15:0] add_ln703_106_fu_4994_p2;
wire   [15:0] add_ln703_107_fu_5000_p2;
wire   [15:0] add_ln703_108_fu_5008_p2;
wire   [15:0] add_ln703_109_fu_5014_p2;
wire   [15:0] add_ln703_110_fu_5022_p2;
wire   [15:0] add_ln703_111_fu_5031_p2;
wire   [15:0] add_ln703_112_fu_5040_p2;
wire   [15:0] add_ln703_113_fu_5049_p2;
wire   [15:0] add_ln703_114_fu_5055_p2;
wire   [15:0] add_ln703_115_fu_5060_p2;
wire   [15:0] add_ln703_116_fu_5068_p2;
wire   [15:0] add_ln703_117_fu_5074_p2;
wire   [15:0] add_ln703_118_fu_5082_p2;
wire   [15:0] add_ln703_119_fu_5091_p2;
wire   [15:0] add_ln703_120_fu_5100_p2;
wire   [15:0] add_ln703_121_fu_5109_p2;
wire   [15:0] add_ln703_122_fu_5118_p2;
wire   [15:0] add_ln703_123_fu_5127_p2;
wire   [15:0] add_ln703_124_fu_5136_p2;
wire   [15:0] add_ln703_125_fu_5145_p2;
wire   [15:0] sext_ln703_3_fu_5160_p1;
wire   [15:0] add_ln703_127_fu_5167_p2;
wire   [15:0] add_ln703_128_fu_5176_p2;
wire   [15:0] add_ln703_129_fu_5182_p2;
reg    grp_fu_428_ce;
reg    grp_fu_430_ce;
reg    grp_fu_431_ce;
reg    grp_fu_432_ce;
reg    grp_fu_433_ce;
reg    grp_fu_435_ce;
reg    grp_fu_436_ce;
reg    grp_fu_437_ce;
reg    grp_fu_438_ce;
reg    grp_fu_439_ce;
reg    grp_fu_440_ce;
reg    grp_fu_441_ce;
reg    grp_fu_442_ce;
reg    grp_fu_443_ce;
reg    grp_fu_444_ce;
reg    grp_fu_445_ce;
reg    grp_fu_446_ce;
reg    grp_fu_447_ce;
reg    grp_fu_448_ce;
reg    grp_fu_449_ce;
reg    grp_fu_451_ce;
reg    grp_fu_452_ce;
reg    grp_fu_453_ce;
reg    grp_fu_454_ce;
reg    grp_fu_455_ce;
reg    grp_fu_456_ce;
reg    grp_fu_457_ce;
reg    grp_fu_458_ce;
reg    grp_fu_459_ce;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U258(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_14_V_read_int_reg),
    .din1(grp_fu_428_p1),
    .ce(grp_fu_428_ce),
    .dout(grp_fu_428_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U259(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_21_V_read_int_reg),
    .din1(grp_fu_430_p1),
    .ce(grp_fu_430_ce),
    .dout(grp_fu_430_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U260(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_13_V_read_int_reg),
    .din1(grp_fu_431_p1),
    .ce(grp_fu_431_ce),
    .dout(grp_fu_431_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U261(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_30_V_read_int_reg),
    .din1(grp_fu_432_p1),
    .ce(grp_fu_432_ce),
    .dout(grp_fu_432_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U262(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_18_V_read_int_reg),
    .din1(grp_fu_433_p1),
    .ce(grp_fu_433_ce),
    .dout(grp_fu_433_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U263(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_0_V_read_int_reg),
    .din1(grp_fu_435_p1),
    .ce(grp_fu_435_ce),
    .dout(grp_fu_435_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U264(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_8_V_read_int_reg),
    .din1(grp_fu_436_p1),
    .ce(grp_fu_436_ce),
    .dout(grp_fu_436_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U265(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_6_V_read_int_reg),
    .din1(grp_fu_437_p1),
    .ce(grp_fu_437_ce),
    .dout(grp_fu_437_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U266(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_11_V_read_int_reg),
    .din1(grp_fu_438_p1),
    .ce(grp_fu_438_ce),
    .dout(grp_fu_438_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U267(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_17_V_read_int_reg),
    .din1(grp_fu_439_p1),
    .ce(grp_fu_439_ce),
    .dout(grp_fu_439_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U268(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_31_V_read_int_reg),
    .din1(grp_fu_440_p1),
    .ce(grp_fu_440_ce),
    .dout(grp_fu_440_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U269(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_25_V_read_int_reg),
    .din1(grp_fu_441_p1),
    .ce(grp_fu_441_ce),
    .dout(grp_fu_441_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U270(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_1_V_read_int_reg),
    .din1(grp_fu_442_p1),
    .ce(grp_fu_442_ce),
    .dout(grp_fu_442_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U271(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_12_V_read_int_reg),
    .din1(grp_fu_443_p1),
    .ce(grp_fu_443_ce),
    .dout(grp_fu_443_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U272(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_4_V_read_int_reg),
    .din1(grp_fu_444_p1),
    .ce(grp_fu_444_ce),
    .dout(grp_fu_444_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U273(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_9_V_read_int_reg),
    .din1(grp_fu_445_p1),
    .ce(grp_fu_445_ce),
    .dout(grp_fu_445_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U274(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_2_V_read_int_reg),
    .din1(grp_fu_446_p1),
    .ce(grp_fu_446_ce),
    .dout(grp_fu_446_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U275(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_23_V_read_int_reg),
    .din1(grp_fu_447_p1),
    .ce(grp_fu_447_ce),
    .dout(grp_fu_447_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U276(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_10_V_read_int_reg),
    .din1(grp_fu_448_p1),
    .ce(grp_fu_448_ce),
    .dout(grp_fu_448_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U277(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_24_V_read_int_reg),
    .din1(grp_fu_449_p1),
    .ce(grp_fu_449_ce),
    .dout(grp_fu_449_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U278(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_20_V_read_int_reg),
    .din1(grp_fu_451_p1),
    .ce(grp_fu_451_ce),
    .dout(grp_fu_451_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U279(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_7_V_read_int_reg),
    .din1(grp_fu_452_p1),
    .ce(grp_fu_452_ce),
    .dout(grp_fu_452_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U280(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_19_V_read_int_reg),
    .din1(grp_fu_453_p1),
    .ce(grp_fu_453_ce),
    .dout(grp_fu_453_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U281(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_5_V_read_int_reg),
    .din1(grp_fu_454_p1),
    .ce(grp_fu_454_ce),
    .dout(grp_fu_454_p2)
);

myproject_mul_16s_10ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_10ns_26_2_0_U282(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_16_V_read_int_reg),
    .din1(grp_fu_455_p1),
    .ce(grp_fu_455_ce),
    .dout(grp_fu_455_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U283(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_15_V_read_int_reg),
    .din1(grp_fu_456_p1),
    .ce(grp_fu_456_ce),
    .dout(grp_fu_456_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U284(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_29_V_read_int_reg),
    .din1(grp_fu_457_p1),
    .ce(grp_fu_457_ce),
    .dout(grp_fu_457_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U285(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_3_V_read_int_reg),
    .din1(grp_fu_458_p1),
    .ce(grp_fu_458_ce),
    .dout(grp_fu_458_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U286(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_26_V_read_int_reg),
    .din1(grp_fu_459_p1),
    .ce(grp_fu_459_ce),
    .dout(grp_fu_459_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_fu_4926_p2;
        ap_return_10_int_reg <= add_ln703_108_fu_5008_p2;
        ap_return_11_int_reg <= add_ln703_109_fu_5014_p2;
        ap_return_12_int_reg <= add_ln703_110_fu_5022_p2;
        ap_return_13_int_reg <= add_ln703_111_fu_5031_p2;
        ap_return_14_int_reg <= add_ln703_112_fu_5040_p2;
        ap_return_15_int_reg <= add_ln703_113_fu_5049_p2;
        ap_return_16_int_reg <= add_ln703_114_fu_5055_p2;
        ap_return_17_int_reg <= add_ln703_115_fu_5060_p2;
        ap_return_18_int_reg <= add_ln703_116_fu_5068_p2;
        ap_return_19_int_reg <= add_ln703_117_fu_5074_p2;
        ap_return_1_int_reg <= add_ln703_99_fu_4935_p2;
        ap_return_20_int_reg <= add_ln703_118_fu_5082_p2;
        ap_return_21_int_reg <= add_ln703_119_fu_5091_p2;
        ap_return_22_int_reg <= add_ln703_120_fu_5100_p2;
        ap_return_23_int_reg <= add_ln703_121_fu_5109_p2;
        ap_return_24_int_reg <= add_ln703_122_fu_5118_p2;
        ap_return_25_int_reg <= add_ln703_123_fu_5127_p2;
        ap_return_26_int_reg <= add_ln703_124_fu_5136_p2;
        ap_return_27_int_reg <= add_ln703_125_fu_5145_p2;
        ap_return_28_int_reg <= sext_ln703_3_fu_5160_p1;
        ap_return_29_int_reg <= add_ln703_127_fu_5167_p2;
        ap_return_2_int_reg <= add_ln703_100_fu_4944_p2;
        ap_return_30_int_reg <= add_ln703_128_fu_5176_p2;
        ap_return_31_int_reg <= add_ln703_129_fu_5182_p2;
        ap_return_3_int_reg <= add_ln703_101_fu_4953_p2;
        ap_return_4_int_reg <= add_ln703_102_fu_4962_p2;
        ap_return_5_int_reg <= add_ln703_103_fu_4971_p2;
        ap_return_6_int_reg <= add_ln703_104_fu_4977_p2;
        ap_return_7_int_reg <= add_ln703_105_fu_4985_p2;
        ap_return_8_int_reg <= add_ln703_106_fu_4994_p2;
        ap_return_9_int_reg <= add_ln703_107_fu_5000_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        tmp_386_reg_5519 <= {{add_ln1118_2_fu_4602_p2[23:10]}};
        tmp_386_reg_5519_pp0_iter1_reg <= tmp_386_reg_5519;
        trunc_ln708_10_reg_5589 <= {{grp_fu_448_p2[24:10]}};
        trunc_ln708_11_reg_5594 <= {{grp_fu_438_p2[25:10]}};
        trunc_ln708_12_reg_5599 <= {{grp_fu_443_p2[24:10]}};
        trunc_ln708_13_reg_5604 <= {{grp_fu_431_p2[24:10]}};
        trunc_ln708_14_reg_5609 <= {{grp_fu_428_p2[24:10]}};
        trunc_ln708_15_reg_5614 <= {{grp_fu_456_p2[24:10]}};
        trunc_ln708_16_reg_5619 <= {{grp_fu_455_p2[25:10]}};
        trunc_ln708_17_reg_5624 <= {{grp_fu_439_p2[25:10]}};
        trunc_ln708_18_reg_5629 <= {{grp_fu_433_p2[24:10]}};
        trunc_ln708_19_reg_5634 <= {{grp_fu_453_p2[25:10]}};
        trunc_ln708_1_reg_5544 <= {{grp_fu_442_p2[24:10]}};
        trunc_ln708_20_reg_5639 <= {{grp_fu_451_p2[24:10]}};
        trunc_ln708_21_reg_5644 <= {{grp_fu_430_p2[24:10]}};
        trunc_ln708_22_reg_5489 <= {{add_ln1118_fu_4502_p2[24:10]}};
        trunc_ln708_22_reg_5489_pp0_iter1_reg <= trunc_ln708_22_reg_5489;
        trunc_ln708_23_reg_5649 <= {{grp_fu_447_p2[24:10]}};
        trunc_ln708_24_reg_5654 <= {{grp_fu_449_p2[24:10]}};
        trunc_ln708_25_reg_5659 <= {{grp_fu_441_p2[24:10]}};
        trunc_ln708_26_reg_5664 <= {{grp_fu_459_p2[24:10]}};
        trunc_ln708_27_reg_5514 <= {{add_ln1118_1_fu_4562_p2[24:10]}};
        trunc_ln708_27_reg_5514_pp0_iter1_reg <= trunc_ln708_27_reg_5514;
        trunc_ln708_29_reg_5669 <= {{grp_fu_457_p2[24:10]}};
        trunc_ln708_2_reg_5549 <= {{grp_fu_446_p2[24:10]}};
        trunc_ln708_30_reg_5674 <= {{grp_fu_432_p2[24:10]}};
        trunc_ln708_31_reg_5679 <= {{grp_fu_440_p2[25:10]}};
        trunc_ln708_3_reg_5554 <= {{grp_fu_458_p2[24:10]}};
        trunc_ln708_4_reg_5559 <= {{grp_fu_444_p2[24:10]}};
        trunc_ln708_5_reg_5564 <= {{grp_fu_454_p2[24:10]}};
        trunc_ln708_6_reg_5569 <= {{grp_fu_437_p2[25:10]}};
        trunc_ln708_7_reg_5574 <= {{grp_fu_452_p2[24:10]}};
        trunc_ln708_8_reg_5579 <= {{grp_fu_436_p2[24:10]}};
        trunc_ln708_9_reg_5584 <= {{grp_fu_445_p2[25:10]}};
        trunc_ln_reg_5539 <= {{grp_fu_435_p2[24:10]}};
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_fu_4926_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = add_ln703_99_fu_4935_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = add_ln703_108_fu_5008_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = add_ln703_109_fu_5014_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = add_ln703_110_fu_5022_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = add_ln703_111_fu_5031_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = add_ln703_112_fu_5040_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = add_ln703_113_fu_5049_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = add_ln703_114_fu_5055_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = add_ln703_115_fu_5060_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = add_ln703_116_fu_5068_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = add_ln703_117_fu_5074_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = add_ln703_100_fu_4944_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = add_ln703_118_fu_5082_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = add_ln703_119_fu_5091_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = add_ln703_120_fu_5100_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = add_ln703_121_fu_5109_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = add_ln703_122_fu_5118_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = add_ln703_123_fu_5127_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = add_ln703_124_fu_5136_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = add_ln703_125_fu_5145_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = sext_ln703_3_fu_5160_p1;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = add_ln703_127_fu_5167_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = add_ln703_101_fu_4953_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = add_ln703_128_fu_5176_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = add_ln703_129_fu_5182_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = add_ln703_102_fu_4962_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = add_ln703_103_fu_4971_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = add_ln703_104_fu_4977_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = add_ln703_105_fu_4985_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = add_ln703_106_fu_4994_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = add_ln703_107_fu_5000_p2;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_428_ce = 1'b1;
    end else begin
        grp_fu_428_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_430_ce = 1'b1;
    end else begin
        grp_fu_430_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_431_ce = 1'b1;
    end else begin
        grp_fu_431_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_432_ce = 1'b1;
    end else begin
        grp_fu_432_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_433_ce = 1'b1;
    end else begin
        grp_fu_433_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_435_ce = 1'b1;
    end else begin
        grp_fu_435_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_436_ce = 1'b1;
    end else begin
        grp_fu_436_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_437_ce = 1'b1;
    end else begin
        grp_fu_437_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_438_ce = 1'b1;
    end else begin
        grp_fu_438_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_439_ce = 1'b1;
    end else begin
        grp_fu_439_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_440_ce = 1'b1;
    end else begin
        grp_fu_440_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_441_ce = 1'b1;
    end else begin
        grp_fu_441_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_442_ce = 1'b1;
    end else begin
        grp_fu_442_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_443_ce = 1'b1;
    end else begin
        grp_fu_443_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_444_ce = 1'b1;
    end else begin
        grp_fu_444_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_445_ce = 1'b1;
    end else begin
        grp_fu_445_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_446_ce = 1'b1;
    end else begin
        grp_fu_446_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_447_ce = 1'b1;
    end else begin
        grp_fu_447_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_448_ce = 1'b1;
    end else begin
        grp_fu_448_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_449_ce = 1'b1;
    end else begin
        grp_fu_449_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_451_ce = 1'b1;
    end else begin
        grp_fu_451_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_452_ce = 1'b1;
    end else begin
        grp_fu_452_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_453_ce = 1'b1;
    end else begin
        grp_fu_453_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_454_ce = 1'b1;
    end else begin
        grp_fu_454_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_455_ce = 1'b1;
    end else begin
        grp_fu_455_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_456_ce = 1'b1;
    end else begin
        grp_fu_456_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_457_ce = 1'b1;
    end else begin
        grp_fu_457_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_458_ce = 1'b1;
    end else begin
        grp_fu_458_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_459_ce = 1'b1;
    end else begin
        grp_fu_459_ce = 1'b0;
    end
end

assign add_ln1118_1_fu_4562_p2 = ((sext_ln1118_29_fu_4558_p1) + (sext_ln1118_28_fu_4546_p1));

assign add_ln1118_2_fu_4602_p2 = ((sext_ln1118_31_fu_4598_p1) + (sext_ln1118_30_fu_4586_p1));

assign add_ln1118_fu_4502_p2 = ((sext_ln1118_23_fu_4498_p1) + (sext_ln1118_22_fu_4486_p1));

assign add_ln703_100_fu_4944_p2 = ((sext_ln708_2_fu_4941_p1) + (16'd176));

assign add_ln703_101_fu_4953_p2 = ((sext_ln708_3_fu_4950_p1) + (16'd64535));

assign add_ln703_102_fu_4962_p2 = ((sext_ln708_4_fu_4959_p1) + (16'd65060));

assign add_ln703_103_fu_4971_p2 = ((sext_ln708_5_fu_4968_p1) + (16'd65037));

assign add_ln703_104_fu_4977_p2 = (trunc_ln708_6_reg_5569 + 16'd1387);

assign add_ln703_105_fu_4985_p2 = ((sext_ln708_6_fu_4982_p1) + (16'd179));

assign add_ln703_106_fu_4994_p2 = ((sext_ln708_7_fu_4991_p1) + (16'd65351));

assign add_ln703_107_fu_5000_p2 = ((trunc_ln708_9_reg_5584) + (16'd64930));

assign add_ln703_108_fu_5008_p2 = ((sext_ln708_8_fu_5005_p1) + (16'd725));

assign add_ln703_109_fu_5014_p2 = ((trunc_ln708_11_reg_5594) + (16'd65311));

assign add_ln703_110_fu_5022_p2 = ((sext_ln708_9_fu_5019_p1) + (16'd419));

assign add_ln703_111_fu_5031_p2 = ((sext_ln708_10_fu_5028_p1) + (16'd64983));

assign add_ln703_112_fu_5040_p2 = ((sext_ln708_11_fu_5037_p1) + (16'd25));

assign add_ln703_113_fu_5049_p2 = ((sext_ln708_12_fu_5046_p1) + (16'd346));

assign add_ln703_114_fu_5055_p2 = (trunc_ln708_16_reg_5619 + 16'd474);

assign add_ln703_115_fu_5060_p2 = ((trunc_ln708_17_reg_5624) + (16'd64364));

assign add_ln703_116_fu_5068_p2 = ((sext_ln708_13_fu_5065_p1) + (16'd65227));

assign add_ln703_117_fu_5074_p2 = (trunc_ln708_19_reg_5634 + 16'd881);

assign add_ln703_118_fu_5082_p2 = ((sext_ln708_14_fu_5079_p1) + (16'd511));

assign add_ln703_119_fu_5091_p2 = ((sext_ln708_15_fu_5088_p1) + (16'd64887));

assign add_ln703_120_fu_5100_p2 = ((sext_ln708_16_fu_5097_p1) + (16'd65275));

assign add_ln703_121_fu_5109_p2 = ((sext_ln708_17_fu_5106_p1) + (16'd664));

assign add_ln703_122_fu_5118_p2 = ((sext_ln708_18_fu_5115_p1) + (16'd513));

assign add_ln703_123_fu_5127_p2 = ((sext_ln708_19_fu_5124_p1) + (16'd833));

assign add_ln703_124_fu_5136_p2 = ((sext_ln708_20_fu_5133_p1) + (16'd332));

assign add_ln703_125_fu_5145_p2 = ((sext_ln708_21_fu_5142_p1) + (16'd65271));

assign add_ln703_126_fu_5154_p2 = ((sext_ln703_fu_5151_p1) + (15'd32312));

assign add_ln703_127_fu_5167_p2 = ((sext_ln708_22_fu_5164_p1) + (16'd423));

assign add_ln703_128_fu_5176_p2 = ((sext_ln708_23_fu_5173_p1) + (16'd399));

assign add_ln703_129_fu_5182_p2 = ((trunc_ln708_31_reg_5679) + (16'd65410));

assign add_ln703_99_fu_4935_p2 = ((sext_ln708_1_fu_4932_p1) + (16'd64428));

assign add_ln703_fu_4926_p2 = ((sext_ln708_fu_4923_p1) + (16'd316));

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign grp_fu_428_p1 = 25'd183;

assign grp_fu_430_p1 = 25'd161;

assign grp_fu_431_p1 = 25'd206;

assign grp_fu_432_p1 = 25'd215;

assign grp_fu_433_p1 = 25'd189;

assign grp_fu_435_p1 = 25'd199;

assign grp_fu_436_p1 = 25'd185;

assign grp_fu_437_p1 = 26'd356;

assign grp_fu_438_p1 = 26'd338;

assign grp_fu_439_p1 = 26'd308;

assign grp_fu_440_p1 = 26'd394;

assign grp_fu_441_p1 = 25'd239;

assign grp_fu_442_p1 = 25'd222;

assign grp_fu_443_p1 = 25'd142;

assign grp_fu_444_p1 = 25'd239;

assign grp_fu_445_p1 = 26'd310;

assign grp_fu_446_p1 = 25'd231;

assign grp_fu_447_p1 = 25'd134;

assign grp_fu_448_p1 = 25'd225;

assign grp_fu_449_p1 = 25'd209;

assign grp_fu_451_p1 = 25'd140;

assign grp_fu_452_p1 = 25'd228;

assign grp_fu_453_p1 = 26'd380;

assign grp_fu_454_p1 = 25'd145;

assign grp_fu_455_p1 = 26'd393;

assign grp_fu_456_p1 = 25'd241;

assign grp_fu_457_p1 = 25'd169;

assign grp_fu_458_p1 = 25'd241;

assign grp_fu_459_p1 = 25'd233;

assign sext_ln1118_22_fu_4486_p0 = data_22_V_read_int_reg;

assign sext_ln1118_22_fu_4486_p1 = sext_ln1118_22_fu_4486_p0;

assign sext_ln1118_23_fu_4498_p1 = (shl_ln_fu_4490_p3);

assign sext_ln1118_28_fu_4546_p1 = (shl_ln1118_1_fu_4538_p3);

assign sext_ln1118_29_fu_4558_p1 = (shl_ln1118_2_fu_4550_p3);

assign sext_ln1118_30_fu_4586_p1 = (shl_ln1118_3_fu_4578_p3);

assign sext_ln1118_31_fu_4598_p1 = (shl_ln1118_4_fu_4590_p3);

assign sext_ln703_3_fu_5160_p1 = (add_ln703_126_fu_5154_p2);

assign sext_ln703_fu_5151_p1 = (tmp_386_reg_5519_pp0_iter1_reg);

assign sext_ln708_10_fu_5028_p1 = (trunc_ln708_13_reg_5604);

assign sext_ln708_11_fu_5037_p1 = (trunc_ln708_14_reg_5609);

assign sext_ln708_12_fu_5046_p1 = (trunc_ln708_15_reg_5614);

assign sext_ln708_13_fu_5065_p1 = (trunc_ln708_18_reg_5629);

assign sext_ln708_14_fu_5079_p1 = (trunc_ln708_20_reg_5639);

assign sext_ln708_15_fu_5088_p1 = (trunc_ln708_21_reg_5644);

assign sext_ln708_16_fu_5097_p1 = (trunc_ln708_22_reg_5489_pp0_iter1_reg);

assign sext_ln708_17_fu_5106_p1 = (trunc_ln708_23_reg_5649);

assign sext_ln708_18_fu_5115_p1 = (trunc_ln708_24_reg_5654);

assign sext_ln708_19_fu_5124_p1 = (trunc_ln708_25_reg_5659);

assign sext_ln708_1_fu_4932_p1 = (trunc_ln708_1_reg_5544);

assign sext_ln708_20_fu_5133_p1 = (trunc_ln708_26_reg_5664);

assign sext_ln708_21_fu_5142_p1 = (trunc_ln708_27_reg_5514_pp0_iter1_reg);

assign sext_ln708_22_fu_5164_p1 = (trunc_ln708_29_reg_5669);

assign sext_ln708_23_fu_5173_p1 = (trunc_ln708_30_reg_5674);

assign sext_ln708_2_fu_4941_p1 = (trunc_ln708_2_reg_5549);

assign sext_ln708_3_fu_4950_p1 = (trunc_ln708_3_reg_5554);

assign sext_ln708_4_fu_4959_p1 = (trunc_ln708_4_reg_5559);

assign sext_ln708_5_fu_4968_p1 = (trunc_ln708_5_reg_5564);

assign sext_ln708_6_fu_4982_p1 = (trunc_ln708_7_reg_5574);

assign sext_ln708_7_fu_4991_p1 = (trunc_ln708_8_reg_5579);

assign sext_ln708_8_fu_5005_p1 = (trunc_ln708_10_reg_5589);

assign sext_ln708_9_fu_5019_p1 = (trunc_ln708_12_reg_5599);

assign sext_ln708_fu_4923_p1 = (trunc_ln_reg_5539);

assign shl_ln1118_1_fu_4538_p3 = {{data_27_V_read_int_reg}, {8'd0}};

assign shl_ln1118_2_fu_4550_p3 = {{data_27_V_read_int_reg}, {6'd0}};

assign shl_ln1118_3_fu_4578_p3 = {{data_28_V_read_int_reg}, {7'd0}};

assign shl_ln1118_4_fu_4590_p3 = {{data_28_V_read_int_reg}, {5'd0}};

assign shl_ln_fu_4490_p1 = data_22_V_read_int_reg;

assign shl_ln_fu_4490_p3 = {{shl_ln_fu_4490_p1}, {8'd0}};

endmodule //normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;

wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [12:0] trunc_ln708_s_reg_362;
reg   [12:0] trunc_ln708_s_reg_362_pp0_iter1_reg;
reg   [14:0] trunc_ln_reg_382;
reg   [14:0] trunc_ln708_1_reg_387;
reg   [14:0] trunc_ln708_2_reg_392;
reg   [14:0] trunc_ln708_3_reg_397;
wire   [8:0] grp_fu_95_p1;
wire    ap_block_pp0_stage0;
wire   [8:0] grp_fu_96_p1;
wire   [8:0] grp_fu_97_p1;
wire   [8:0] grp_fu_98_p1;
wire   [24:0] grp_fu_98_p2;
wire   [24:0] grp_fu_96_p2;
wire   [24:0] grp_fu_97_p2;
wire   [24:0] grp_fu_95_p2;
wire   [15:0] sext_ln708_fu_278_p1;
wire   [13:0] sext_ln703_fu_287_p1;
wire   [13:0] add_ln703_1_fu_290_p2;
wire   [15:0] sext_ln708_1_fu_300_p1;
wire   [15:0] sext_ln708_2_fu_309_p1;
wire   [15:0] sext_ln708_3_fu_318_p1;
wire   [15:0] add_ln703_fu_281_p2;
wire   [15:0] sext_ln703_1_fu_296_p1;
wire   [15:0] add_ln703_2_fu_303_p2;
wire   [15:0] add_ln703_3_fu_312_p2;
wire   [15:0] add_ln703_4_fu_321_p2;
reg    grp_fu_95_ce;
reg    grp_fu_96_ce;
reg    grp_fu_97_ce;
reg    grp_fu_98_ce;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U513(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_4_V_read_int_reg),
    .din1(grp_fu_95_p1),
    .ce(grp_fu_95_ce),
    .dout(grp_fu_95_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U514(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_2_V_read_int_reg),
    .din1(grp_fu_96_p1),
    .ce(grp_fu_96_ce),
    .dout(grp_fu_96_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U515(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_3_V_read_int_reg),
    .din1(grp_fu_97_p1),
    .ce(grp_fu_97_ce),
    .dout(grp_fu_97_p2)
);

myproject_mul_16s_9ns_25_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 25 ))
myproject_mul_16s_9ns_25_2_0_U516(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_0_V_read_int_reg),
    .din1(grp_fu_98_p1),
    .ce(grp_fu_98_ce),
    .dout(grp_fu_98_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_fu_281_p2;
        ap_return_1_int_reg <= sext_ln703_1_fu_296_p1;
        ap_return_2_int_reg <= add_ln703_2_fu_303_p2;
        ap_return_3_int_reg <= add_ln703_3_fu_312_p2;
        ap_return_4_int_reg <= add_ln703_4_fu_321_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        trunc_ln708_1_reg_387 <= {{grp_fu_96_p2[24:10]}};
        trunc_ln708_2_reg_392 <= {{grp_fu_97_p2[24:10]}};
        trunc_ln708_3_reg_397 <= {{grp_fu_95_p2[24:10]}};
        trunc_ln708_s_reg_362 <= {{data_1_V_read_int_reg[15:3]}};
        trunc_ln708_s_reg_362_pp0_iter1_reg <= trunc_ln708_s_reg_362;
        trunc_ln_reg_382 <= {{grp_fu_98_p2[24:10]}};
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_fu_281_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = sext_ln703_1_fu_296_p1;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = add_ln703_2_fu_303_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = add_ln703_3_fu_312_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = add_ln703_4_fu_321_p2;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_95_ce = 1'b1;
    end else begin
        grp_fu_95_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_96_ce = 1'b1;
    end else begin
        grp_fu_96_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_97_ce = 1'b1;
    end else begin
        grp_fu_97_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        grp_fu_98_ce = 1'b1;
    end else begin
        grp_fu_98_ce = 1'b0;
    end
end

assign add_ln703_1_fu_290_p2 = ((sext_ln703_fu_287_p1) + (14'd15560));

assign add_ln703_2_fu_303_p2 = ((sext_ln708_1_fu_300_p1) + (16'd64405));

assign add_ln703_3_fu_312_p2 = ((sext_ln708_2_fu_309_p1) + (16'd64656));

assign add_ln703_4_fu_321_p2 = ((sext_ln708_3_fu_318_p1) + (16'd65325));

assign add_ln703_fu_281_p2 = ((sext_ln708_fu_278_p1) + (16'd64860));

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign grp_fu_95_p1 = 25'd162;

assign grp_fu_96_p1 = 25'd239;

assign grp_fu_97_p1 = 25'd221;

assign grp_fu_98_p1 = 25'd174;

assign sext_ln703_1_fu_296_p1 = (add_ln703_1_fu_290_p2);

assign sext_ln703_fu_287_p1 = (trunc_ln708_s_reg_362_pp0_iter1_reg);

assign sext_ln708_1_fu_300_p1 = (trunc_ln708_1_reg_387);

assign sext_ln708_2_fu_309_p1 = (trunc_ln708_2_reg_392);

assign sext_ln708_3_fu_318_p1 = (trunc_ln708_3_reg_397);

assign sext_ln708_fu_278_p1 = (trunc_ln_reg_382);

endmodule //normalize_ap_fixed_ap_fixed_config16_0_0_0_0_0_0_0_0_0_0
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module relu_max_ap_fixed_ap_fixed_1_relu1_config13_s (
        ap_ready,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31
);


output   ap_ready;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;

wire   [0:0] tmp_290_fu_302_p3;
wire   [0:0] xor_ln1495_fu_310_p2;
wire   [10:0] tmp_291_fu_316_p3;
wire   [0:0] tmp_289_fu_288_p3;
wire   [0:0] icmp_ln1494_fu_296_p2;
wire   [0:0] or_ln1495_fu_328_p2;
wire   [15:0] zext_ln1495_fu_324_p1;
wire   [0:0] tmp_293_fu_356_p3;
wire   [0:0] xor_ln1495_95_fu_364_p2;
wire   [10:0] tmp_294_fu_370_p3;
wire   [0:0] tmp_292_fu_342_p3;
wire   [0:0] icmp_ln1494_1_fu_350_p2;
wire   [0:0] or_ln1495_95_fu_382_p2;
wire   [15:0] zext_ln1495_95_fu_378_p1;
wire   [0:0] tmp_296_fu_410_p3;
wire   [0:0] xor_ln1495_96_fu_418_p2;
wire   [10:0] tmp_297_fu_424_p3;
wire   [0:0] tmp_295_fu_396_p3;
wire   [0:0] icmp_ln1494_2_fu_404_p2;
wire   [0:0] or_ln1495_96_fu_436_p2;
wire   [15:0] zext_ln1495_96_fu_432_p1;
wire   [0:0] tmp_299_fu_464_p3;
wire   [0:0] xor_ln1495_97_fu_472_p2;
wire   [10:0] tmp_300_fu_478_p3;
wire   [0:0] tmp_298_fu_450_p3;
wire   [0:0] icmp_ln1494_3_fu_458_p2;
wire   [0:0] or_ln1495_97_fu_490_p2;
wire   [15:0] zext_ln1495_97_fu_486_p1;
wire   [0:0] tmp_302_fu_518_p3;
wire   [0:0] xor_ln1495_98_fu_526_p2;
wire   [10:0] tmp_303_fu_532_p3;
wire   [0:0] tmp_301_fu_504_p3;
wire   [0:0] icmp_ln1494_4_fu_512_p2;
wire   [0:0] or_ln1495_98_fu_544_p2;
wire   [15:0] zext_ln1495_98_fu_540_p1;
wire   [0:0] tmp_305_fu_572_p3;
wire   [0:0] xor_ln1495_99_fu_580_p2;
wire   [10:0] tmp_306_fu_586_p3;
wire   [0:0] tmp_304_fu_558_p3;
wire   [0:0] icmp_ln1494_5_fu_566_p2;
wire   [0:0] or_ln1495_99_fu_598_p2;
wire   [15:0] zext_ln1495_99_fu_594_p1;
wire   [0:0] tmp_308_fu_626_p3;
wire   [0:0] xor_ln1495_100_fu_634_p2;
wire   [10:0] tmp_309_fu_640_p3;
wire   [0:0] tmp_307_fu_612_p3;
wire   [0:0] icmp_ln1494_6_fu_620_p2;
wire   [0:0] or_ln1495_100_fu_652_p2;
wire   [15:0] zext_ln1495_100_fu_648_p1;
wire   [0:0] tmp_311_fu_680_p3;
wire   [0:0] xor_ln1495_101_fu_688_p2;
wire   [10:0] tmp_312_fu_694_p3;
wire   [0:0] tmp_310_fu_666_p3;
wire   [0:0] icmp_ln1494_7_fu_674_p2;
wire   [0:0] or_ln1495_101_fu_706_p2;
wire   [15:0] zext_ln1495_101_fu_702_p1;
wire   [0:0] tmp_314_fu_734_p3;
wire   [0:0] xor_ln1495_102_fu_742_p2;
wire   [10:0] tmp_315_fu_748_p3;
wire   [0:0] tmp_313_fu_720_p3;
wire   [0:0] icmp_ln1494_8_fu_728_p2;
wire   [0:0] or_ln1495_102_fu_760_p2;
wire   [15:0] zext_ln1495_102_fu_756_p1;
wire   [0:0] tmp_317_fu_788_p3;
wire   [0:0] xor_ln1495_103_fu_796_p2;
wire   [10:0] tmp_318_fu_802_p3;
wire   [0:0] tmp_316_fu_774_p3;
wire   [0:0] icmp_ln1494_9_fu_782_p2;
wire   [0:0] or_ln1495_103_fu_814_p2;
wire   [15:0] zext_ln1495_103_fu_810_p1;
wire   [0:0] tmp_320_fu_842_p3;
wire   [0:0] xor_ln1495_104_fu_850_p2;
wire   [10:0] tmp_321_fu_856_p3;
wire   [0:0] tmp_319_fu_828_p3;
wire   [0:0] icmp_ln1494_10_fu_836_p2;
wire   [0:0] or_ln1495_104_fu_868_p2;
wire   [15:0] zext_ln1495_104_fu_864_p1;
wire   [0:0] tmp_323_fu_896_p3;
wire   [0:0] xor_ln1495_105_fu_904_p2;
wire   [10:0] tmp_324_fu_910_p3;
wire   [0:0] tmp_322_fu_882_p3;
wire   [0:0] icmp_ln1494_11_fu_890_p2;
wire   [0:0] or_ln1495_105_fu_922_p2;
wire   [15:0] zext_ln1495_105_fu_918_p1;
wire   [0:0] tmp_326_fu_950_p3;
wire   [0:0] xor_ln1495_106_fu_958_p2;
wire   [10:0] tmp_327_fu_964_p3;
wire   [0:0] tmp_325_fu_936_p3;
wire   [0:0] icmp_ln1494_12_fu_944_p2;
wire   [0:0] or_ln1495_106_fu_976_p2;
wire   [15:0] zext_ln1495_106_fu_972_p1;
wire   [0:0] tmp_329_fu_1004_p3;
wire   [0:0] xor_ln1495_107_fu_1012_p2;
wire   [10:0] tmp_330_fu_1018_p3;
wire   [0:0] tmp_328_fu_990_p3;
wire   [0:0] icmp_ln1494_13_fu_998_p2;
wire   [0:0] or_ln1495_107_fu_1030_p2;
wire   [15:0] zext_ln1495_107_fu_1026_p1;
wire   [0:0] tmp_332_fu_1058_p3;
wire   [0:0] xor_ln1495_108_fu_1066_p2;
wire   [10:0] tmp_333_fu_1072_p3;
wire   [0:0] tmp_331_fu_1044_p3;
wire   [0:0] icmp_ln1494_14_fu_1052_p2;
wire   [0:0] or_ln1495_108_fu_1084_p2;
wire   [15:0] zext_ln1495_108_fu_1080_p1;
wire   [0:0] tmp_335_fu_1112_p3;
wire   [0:0] xor_ln1495_109_fu_1120_p2;
wire   [10:0] tmp_336_fu_1126_p3;
wire   [0:0] tmp_334_fu_1098_p3;
wire   [0:0] icmp_ln1494_15_fu_1106_p2;
wire   [0:0] or_ln1495_109_fu_1138_p2;
wire   [15:0] zext_ln1495_109_fu_1134_p1;
wire   [0:0] tmp_338_fu_1166_p3;
wire   [0:0] xor_ln1495_110_fu_1174_p2;
wire   [10:0] tmp_339_fu_1180_p3;
wire   [0:0] tmp_337_fu_1152_p3;
wire   [0:0] icmp_ln1494_16_fu_1160_p2;
wire   [0:0] or_ln1495_110_fu_1192_p2;
wire   [15:0] zext_ln1495_110_fu_1188_p1;
wire   [0:0] tmp_341_fu_1220_p3;
wire   [0:0] xor_ln1495_111_fu_1228_p2;
wire   [10:0] tmp_342_fu_1234_p3;
wire   [0:0] tmp_340_fu_1206_p3;
wire   [0:0] icmp_ln1494_17_fu_1214_p2;
wire   [0:0] or_ln1495_111_fu_1246_p2;
wire   [15:0] zext_ln1495_111_fu_1242_p1;
wire   [0:0] tmp_344_fu_1274_p3;
wire   [0:0] xor_ln1495_112_fu_1282_p2;
wire   [10:0] tmp_345_fu_1288_p3;
wire   [0:0] tmp_343_fu_1260_p3;
wire   [0:0] icmp_ln1494_18_fu_1268_p2;
wire   [0:0] or_ln1495_112_fu_1300_p2;
wire   [15:0] zext_ln1495_112_fu_1296_p1;
wire   [0:0] tmp_347_fu_1328_p3;
wire   [0:0] xor_ln1495_113_fu_1336_p2;
wire   [10:0] tmp_348_fu_1342_p3;
wire   [0:0] tmp_346_fu_1314_p3;
wire   [0:0] icmp_ln1494_19_fu_1322_p2;
wire   [0:0] or_ln1495_113_fu_1354_p2;
wire   [15:0] zext_ln1495_113_fu_1350_p1;
wire   [0:0] tmp_350_fu_1382_p3;
wire   [0:0] xor_ln1495_114_fu_1390_p2;
wire   [10:0] tmp_351_fu_1396_p3;
wire   [0:0] tmp_349_fu_1368_p3;
wire   [0:0] icmp_ln1494_20_fu_1376_p2;
wire   [0:0] or_ln1495_114_fu_1408_p2;
wire   [15:0] zext_ln1495_114_fu_1404_p1;
wire   [0:0] tmp_353_fu_1436_p3;
wire   [0:0] xor_ln1495_115_fu_1444_p2;
wire   [10:0] tmp_354_fu_1450_p3;
wire   [0:0] tmp_352_fu_1422_p3;
wire   [0:0] icmp_ln1494_21_fu_1430_p2;
wire   [0:0] or_ln1495_115_fu_1462_p2;
wire   [15:0] zext_ln1495_115_fu_1458_p1;
wire   [0:0] tmp_356_fu_1490_p3;
wire   [0:0] xor_ln1495_116_fu_1498_p2;
wire   [10:0] tmp_357_fu_1504_p3;
wire   [0:0] tmp_355_fu_1476_p3;
wire   [0:0] icmp_ln1494_22_fu_1484_p2;
wire   [0:0] or_ln1495_116_fu_1516_p2;
wire   [15:0] zext_ln1495_116_fu_1512_p1;
wire   [0:0] tmp_359_fu_1544_p3;
wire   [0:0] xor_ln1495_117_fu_1552_p2;
wire   [10:0] tmp_360_fu_1558_p3;
wire   [0:0] tmp_358_fu_1530_p3;
wire   [0:0] icmp_ln1494_23_fu_1538_p2;
wire   [0:0] or_ln1495_117_fu_1570_p2;
wire   [15:0] zext_ln1495_117_fu_1566_p1;
wire   [0:0] tmp_362_fu_1598_p3;
wire   [0:0] xor_ln1495_118_fu_1606_p2;
wire   [10:0] tmp_363_fu_1612_p3;
wire   [0:0] tmp_361_fu_1584_p3;
wire   [0:0] icmp_ln1494_24_fu_1592_p2;
wire   [0:0] or_ln1495_118_fu_1624_p2;
wire   [15:0] zext_ln1495_118_fu_1620_p1;
wire   [0:0] tmp_365_fu_1652_p3;
wire   [0:0] xor_ln1495_119_fu_1660_p2;
wire   [10:0] tmp_366_fu_1666_p3;
wire   [0:0] tmp_364_fu_1638_p3;
wire   [0:0] icmp_ln1494_25_fu_1646_p2;
wire   [0:0] or_ln1495_119_fu_1678_p2;
wire   [15:0] zext_ln1495_119_fu_1674_p1;
wire   [0:0] tmp_368_fu_1706_p3;
wire   [0:0] xor_ln1495_120_fu_1714_p2;
wire   [10:0] tmp_369_fu_1720_p3;
wire   [0:0] tmp_367_fu_1692_p3;
wire   [0:0] icmp_ln1494_26_fu_1700_p2;
wire   [0:0] or_ln1495_120_fu_1732_p2;
wire   [15:0] zext_ln1495_120_fu_1728_p1;
wire   [0:0] tmp_371_fu_1760_p3;
wire   [0:0] xor_ln1495_121_fu_1768_p2;
wire   [10:0] tmp_372_fu_1774_p3;
wire   [0:0] tmp_370_fu_1746_p3;
wire   [0:0] icmp_ln1494_27_fu_1754_p2;
wire   [0:0] or_ln1495_121_fu_1786_p2;
wire   [15:0] zext_ln1495_121_fu_1782_p1;
wire   [0:0] tmp_374_fu_1814_p3;
wire   [0:0] xor_ln1495_122_fu_1822_p2;
wire   [10:0] tmp_375_fu_1828_p3;
wire   [0:0] tmp_373_fu_1800_p3;
wire   [0:0] icmp_ln1494_28_fu_1808_p2;
wire   [0:0] or_ln1495_122_fu_1840_p2;
wire   [15:0] zext_ln1495_122_fu_1836_p1;
wire   [0:0] tmp_377_fu_1868_p3;
wire   [0:0] xor_ln1495_123_fu_1876_p2;
wire   [10:0] tmp_378_fu_1882_p3;
wire   [0:0] tmp_376_fu_1854_p3;
wire   [0:0] icmp_ln1494_29_fu_1862_p2;
wire   [0:0] or_ln1495_123_fu_1894_p2;
wire   [15:0] zext_ln1495_123_fu_1890_p1;
wire   [0:0] tmp_380_fu_1922_p3;
wire   [0:0] xor_ln1495_124_fu_1930_p2;
wire   [10:0] tmp_381_fu_1936_p3;
wire   [0:0] tmp_379_fu_1908_p3;
wire   [0:0] icmp_ln1494_30_fu_1916_p2;
wire   [0:0] or_ln1495_124_fu_1948_p2;
wire   [15:0] zext_ln1495_124_fu_1944_p1;
wire   [0:0] tmp_383_fu_1976_p3;
wire   [0:0] xor_ln1495_125_fu_1984_p2;
wire   [10:0] tmp_384_fu_1990_p3;
wire   [0:0] tmp_382_fu_1962_p3;
wire   [0:0] icmp_ln1494_31_fu_1970_p2;
wire   [0:0] or_ln1495_125_fu_2002_p2;
wire   [15:0] zext_ln1495_125_fu_1998_p1;
wire   [15:0] select_ln1495_fu_334_p3;
wire   [15:0] select_ln1495_95_fu_388_p3;
wire   [15:0] select_ln1495_96_fu_442_p3;
wire   [15:0] select_ln1495_97_fu_496_p3;
wire   [15:0] select_ln1495_98_fu_550_p3;
wire   [15:0] select_ln1495_99_fu_604_p3;
wire   [15:0] select_ln1495_100_fu_658_p3;
wire   [15:0] select_ln1495_101_fu_712_p3;
wire   [15:0] select_ln1495_102_fu_766_p3;
wire   [15:0] select_ln1495_103_fu_820_p3;
wire   [15:0] select_ln1495_104_fu_874_p3;
wire   [15:0] select_ln1495_105_fu_928_p3;
wire   [15:0] select_ln1495_106_fu_982_p3;
wire   [15:0] select_ln1495_107_fu_1036_p3;
wire   [15:0] select_ln1495_108_fu_1090_p3;
wire   [15:0] select_ln1495_109_fu_1144_p3;
wire   [15:0] select_ln1495_110_fu_1198_p3;
wire   [15:0] select_ln1495_111_fu_1252_p3;
wire   [15:0] select_ln1495_112_fu_1306_p3;
wire   [15:0] select_ln1495_113_fu_1360_p3;
wire   [15:0] select_ln1495_114_fu_1414_p3;
wire   [15:0] select_ln1495_115_fu_1468_p3;
wire   [15:0] select_ln1495_116_fu_1522_p3;
wire   [15:0] select_ln1495_117_fu_1576_p3;
wire   [15:0] select_ln1495_118_fu_1630_p3;
wire   [15:0] select_ln1495_119_fu_1684_p3;
wire   [15:0] select_ln1495_120_fu_1738_p3;
wire   [15:0] select_ln1495_121_fu_1792_p3;
wire   [15:0] select_ln1495_122_fu_1846_p3;
wire   [15:0] select_ln1495_123_fu_1900_p3;
wire   [15:0] select_ln1495_124_fu_1954_p3;
wire   [15:0] select_ln1495_125_fu_2008_p3;

assign ap_ready = 1'b1;

assign ap_return_0 = select_ln1495_fu_334_p3;

assign ap_return_1 = select_ln1495_95_fu_388_p3;

assign ap_return_10 = select_ln1495_104_fu_874_p3;

assign ap_return_11 = select_ln1495_105_fu_928_p3;

assign ap_return_12 = select_ln1495_106_fu_982_p3;

assign ap_return_13 = select_ln1495_107_fu_1036_p3;

assign ap_return_14 = select_ln1495_108_fu_1090_p3;

assign ap_return_15 = select_ln1495_109_fu_1144_p3;

assign ap_return_16 = select_ln1495_110_fu_1198_p3;

assign ap_return_17 = select_ln1495_111_fu_1252_p3;

assign ap_return_18 = select_ln1495_112_fu_1306_p3;

assign ap_return_19 = select_ln1495_113_fu_1360_p3;

assign ap_return_2 = select_ln1495_96_fu_442_p3;

assign ap_return_20 = select_ln1495_114_fu_1414_p3;

assign ap_return_21 = select_ln1495_115_fu_1468_p3;

assign ap_return_22 = select_ln1495_116_fu_1522_p3;

assign ap_return_23 = select_ln1495_117_fu_1576_p3;

assign ap_return_24 = select_ln1495_118_fu_1630_p3;

assign ap_return_25 = select_ln1495_119_fu_1684_p3;

assign ap_return_26 = select_ln1495_120_fu_1738_p3;

assign ap_return_27 = select_ln1495_121_fu_1792_p3;

assign ap_return_28 = select_ln1495_122_fu_1846_p3;

assign ap_return_29 = select_ln1495_123_fu_1900_p3;

assign ap_return_3 = select_ln1495_97_fu_496_p3;

assign ap_return_30 = select_ln1495_124_fu_1954_p3;

assign ap_return_31 = select_ln1495_125_fu_2008_p3;

assign ap_return_4 = select_ln1495_98_fu_550_p3;

assign ap_return_5 = select_ln1495_99_fu_604_p3;

assign ap_return_6 = select_ln1495_100_fu_658_p3;

assign ap_return_7 = select_ln1495_101_fu_712_p3;

assign ap_return_8 = select_ln1495_102_fu_766_p3;

assign ap_return_9 = select_ln1495_103_fu_820_p3;

assign icmp_ln1494_10_fu_836_p2 = (((data_10_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_11_fu_890_p2 = (((data_11_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_12_fu_944_p2 = (((data_12_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_13_fu_998_p2 = (((data_13_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_14_fu_1052_p2 = (((data_14_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_15_fu_1106_p2 = (((data_15_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_16_fu_1160_p2 = (((data_16_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_17_fu_1214_p2 = (((data_17_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_18_fu_1268_p2 = (((data_18_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_19_fu_1322_p2 = (((data_19_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_1_fu_350_p2 = (((data_1_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_20_fu_1376_p2 = (((data_20_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_21_fu_1430_p2 = (((data_21_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_22_fu_1484_p2 = (((data_22_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_23_fu_1538_p2 = (((data_23_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_24_fu_1592_p2 = (((data_24_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_25_fu_1646_p2 = (((data_25_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_26_fu_1700_p2 = (((data_26_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_27_fu_1754_p2 = (((data_27_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_28_fu_1808_p2 = (((data_28_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_29_fu_1862_p2 = (((data_29_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_2_fu_404_p2 = (((data_2_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_30_fu_1916_p2 = (((data_30_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_31_fu_1970_p2 = (((data_31_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_3_fu_458_p2 = (((data_3_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_4_fu_512_p2 = (((data_4_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_5_fu_566_p2 = (((data_5_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_6_fu_620_p2 = (((data_6_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_7_fu_674_p2 = (((data_7_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_8_fu_728_p2 = (((data_8_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_9_fu_782_p2 = (((data_9_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_fu_296_p2 = (((data_0_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign or_ln1495_100_fu_652_p2 = (tmp_307_fu_612_p3 | icmp_ln1494_6_fu_620_p2);

assign or_ln1495_101_fu_706_p2 = (tmp_310_fu_666_p3 | icmp_ln1494_7_fu_674_p2);

assign or_ln1495_102_fu_760_p2 = (tmp_313_fu_720_p3 | icmp_ln1494_8_fu_728_p2);

assign or_ln1495_103_fu_814_p2 = (tmp_316_fu_774_p3 | icmp_ln1494_9_fu_782_p2);

assign or_ln1495_104_fu_868_p2 = (tmp_319_fu_828_p3 | icmp_ln1494_10_fu_836_p2);

assign or_ln1495_105_fu_922_p2 = (tmp_322_fu_882_p3 | icmp_ln1494_11_fu_890_p2);

assign or_ln1495_106_fu_976_p2 = (tmp_325_fu_936_p3 | icmp_ln1494_12_fu_944_p2);

assign or_ln1495_107_fu_1030_p2 = (tmp_328_fu_990_p3 | icmp_ln1494_13_fu_998_p2);

assign or_ln1495_108_fu_1084_p2 = (tmp_331_fu_1044_p3 | icmp_ln1494_14_fu_1052_p2);

assign or_ln1495_109_fu_1138_p2 = (tmp_334_fu_1098_p3 | icmp_ln1494_15_fu_1106_p2);

assign or_ln1495_110_fu_1192_p2 = (tmp_337_fu_1152_p3 | icmp_ln1494_16_fu_1160_p2);

assign or_ln1495_111_fu_1246_p2 = (tmp_340_fu_1206_p3 | icmp_ln1494_17_fu_1214_p2);

assign or_ln1495_112_fu_1300_p2 = (tmp_343_fu_1260_p3 | icmp_ln1494_18_fu_1268_p2);

assign or_ln1495_113_fu_1354_p2 = (tmp_346_fu_1314_p3 | icmp_ln1494_19_fu_1322_p2);

assign or_ln1495_114_fu_1408_p2 = (tmp_349_fu_1368_p3 | icmp_ln1494_20_fu_1376_p2);

assign or_ln1495_115_fu_1462_p2 = (tmp_352_fu_1422_p3 | icmp_ln1494_21_fu_1430_p2);

assign or_ln1495_116_fu_1516_p2 = (tmp_355_fu_1476_p3 | icmp_ln1494_22_fu_1484_p2);

assign or_ln1495_117_fu_1570_p2 = (tmp_358_fu_1530_p3 | icmp_ln1494_23_fu_1538_p2);

assign or_ln1495_118_fu_1624_p2 = (tmp_361_fu_1584_p3 | icmp_ln1494_24_fu_1592_p2);

assign or_ln1495_119_fu_1678_p2 = (tmp_364_fu_1638_p3 | icmp_ln1494_25_fu_1646_p2);

assign or_ln1495_120_fu_1732_p2 = (tmp_367_fu_1692_p3 | icmp_ln1494_26_fu_1700_p2);

assign or_ln1495_121_fu_1786_p2 = (tmp_370_fu_1746_p3 | icmp_ln1494_27_fu_1754_p2);

assign or_ln1495_122_fu_1840_p2 = (tmp_373_fu_1800_p3 | icmp_ln1494_28_fu_1808_p2);

assign or_ln1495_123_fu_1894_p2 = (tmp_376_fu_1854_p3 | icmp_ln1494_29_fu_1862_p2);

assign or_ln1495_124_fu_1948_p2 = (tmp_379_fu_1908_p3 | icmp_ln1494_30_fu_1916_p2);

assign or_ln1495_125_fu_2002_p2 = (tmp_382_fu_1962_p3 | icmp_ln1494_31_fu_1970_p2);

assign or_ln1495_95_fu_382_p2 = (tmp_292_fu_342_p3 | icmp_ln1494_1_fu_350_p2);

assign or_ln1495_96_fu_436_p2 = (tmp_295_fu_396_p3 | icmp_ln1494_2_fu_404_p2);

assign or_ln1495_97_fu_490_p2 = (tmp_298_fu_450_p3 | icmp_ln1494_3_fu_458_p2);

assign or_ln1495_98_fu_544_p2 = (tmp_301_fu_504_p3 | icmp_ln1494_4_fu_512_p2);

assign or_ln1495_99_fu_598_p2 = (tmp_304_fu_558_p3 | icmp_ln1494_5_fu_566_p2);

assign or_ln1495_fu_328_p2 = (tmp_289_fu_288_p3 | icmp_ln1494_fu_296_p2);

assign select_ln1495_100_fu_658_p3 = ((or_ln1495_100_fu_652_p2[0:0] == 1'b1) ? zext_ln1495_100_fu_648_p1 : data_6_V_read);

assign select_ln1495_101_fu_712_p3 = ((or_ln1495_101_fu_706_p2[0:0] == 1'b1) ? zext_ln1495_101_fu_702_p1 : data_7_V_read);

assign select_ln1495_102_fu_766_p3 = ((or_ln1495_102_fu_760_p2[0:0] == 1'b1) ? zext_ln1495_102_fu_756_p1 : data_8_V_read);

assign select_ln1495_103_fu_820_p3 = ((or_ln1495_103_fu_814_p2[0:0] == 1'b1) ? zext_ln1495_103_fu_810_p1 : data_9_V_read);

assign select_ln1495_104_fu_874_p3 = ((or_ln1495_104_fu_868_p2[0:0] == 1'b1) ? zext_ln1495_104_fu_864_p1 : data_10_V_read);

assign select_ln1495_105_fu_928_p3 = ((or_ln1495_105_fu_922_p2[0:0] == 1'b1) ? zext_ln1495_105_fu_918_p1 : data_11_V_read);

assign select_ln1495_106_fu_982_p3 = ((or_ln1495_106_fu_976_p2[0:0] == 1'b1) ? zext_ln1495_106_fu_972_p1 : data_12_V_read);

assign select_ln1495_107_fu_1036_p3 = ((or_ln1495_107_fu_1030_p2[0:0] == 1'b1) ? zext_ln1495_107_fu_1026_p1 : data_13_V_read);

assign select_ln1495_108_fu_1090_p3 = ((or_ln1495_108_fu_1084_p2[0:0] == 1'b1) ? zext_ln1495_108_fu_1080_p1 : data_14_V_read);

assign select_ln1495_109_fu_1144_p3 = ((or_ln1495_109_fu_1138_p2[0:0] == 1'b1) ? zext_ln1495_109_fu_1134_p1 : data_15_V_read);

assign select_ln1495_110_fu_1198_p3 = ((or_ln1495_110_fu_1192_p2[0:0] == 1'b1) ? zext_ln1495_110_fu_1188_p1 : data_16_V_read);

assign select_ln1495_111_fu_1252_p3 = ((or_ln1495_111_fu_1246_p2[0:0] == 1'b1) ? zext_ln1495_111_fu_1242_p1 : data_17_V_read);

assign select_ln1495_112_fu_1306_p3 = ((or_ln1495_112_fu_1300_p2[0:0] == 1'b1) ? zext_ln1495_112_fu_1296_p1 : data_18_V_read);

assign select_ln1495_113_fu_1360_p3 = ((or_ln1495_113_fu_1354_p2[0:0] == 1'b1) ? zext_ln1495_113_fu_1350_p1 : data_19_V_read);

assign select_ln1495_114_fu_1414_p3 = ((or_ln1495_114_fu_1408_p2[0:0] == 1'b1) ? zext_ln1495_114_fu_1404_p1 : data_20_V_read);

assign select_ln1495_115_fu_1468_p3 = ((or_ln1495_115_fu_1462_p2[0:0] == 1'b1) ? zext_ln1495_115_fu_1458_p1 : data_21_V_read);

assign select_ln1495_116_fu_1522_p3 = ((or_ln1495_116_fu_1516_p2[0:0] == 1'b1) ? zext_ln1495_116_fu_1512_p1 : data_22_V_read);

assign select_ln1495_117_fu_1576_p3 = ((or_ln1495_117_fu_1570_p2[0:0] == 1'b1) ? zext_ln1495_117_fu_1566_p1 : data_23_V_read);

assign select_ln1495_118_fu_1630_p3 = ((or_ln1495_118_fu_1624_p2[0:0] == 1'b1) ? zext_ln1495_118_fu_1620_p1 : data_24_V_read);

assign select_ln1495_119_fu_1684_p3 = ((or_ln1495_119_fu_1678_p2[0:0] == 1'b1) ? zext_ln1495_119_fu_1674_p1 : data_25_V_read);

assign select_ln1495_120_fu_1738_p3 = ((or_ln1495_120_fu_1732_p2[0:0] == 1'b1) ? zext_ln1495_120_fu_1728_p1 : data_26_V_read);

assign select_ln1495_121_fu_1792_p3 = ((or_ln1495_121_fu_1786_p2[0:0] == 1'b1) ? zext_ln1495_121_fu_1782_p1 : data_27_V_read);

assign select_ln1495_122_fu_1846_p3 = ((or_ln1495_122_fu_1840_p2[0:0] == 1'b1) ? zext_ln1495_122_fu_1836_p1 : data_28_V_read);

assign select_ln1495_123_fu_1900_p3 = ((or_ln1495_123_fu_1894_p2[0:0] == 1'b1) ? zext_ln1495_123_fu_1890_p1 : data_29_V_read);

assign select_ln1495_124_fu_1954_p3 = ((or_ln1495_124_fu_1948_p2[0:0] == 1'b1) ? zext_ln1495_124_fu_1944_p1 : data_30_V_read);

assign select_ln1495_125_fu_2008_p3 = ((or_ln1495_125_fu_2002_p2[0:0] == 1'b1) ? zext_ln1495_125_fu_1998_p1 : data_31_V_read);

assign select_ln1495_95_fu_388_p3 = ((or_ln1495_95_fu_382_p2[0:0] == 1'b1) ? zext_ln1495_95_fu_378_p1 : data_1_V_read);

assign select_ln1495_96_fu_442_p3 = ((or_ln1495_96_fu_436_p2[0:0] == 1'b1) ? zext_ln1495_96_fu_432_p1 : data_2_V_read);

assign select_ln1495_97_fu_496_p3 = ((or_ln1495_97_fu_490_p2[0:0] == 1'b1) ? zext_ln1495_97_fu_486_p1 : data_3_V_read);

assign select_ln1495_98_fu_550_p3 = ((or_ln1495_98_fu_544_p2[0:0] == 1'b1) ? zext_ln1495_98_fu_540_p1 : data_4_V_read);

assign select_ln1495_99_fu_604_p3 = ((or_ln1495_99_fu_598_p2[0:0] == 1'b1) ? zext_ln1495_99_fu_594_p1 : data_5_V_read);

assign select_ln1495_fu_334_p3 = ((or_ln1495_fu_328_p2[0:0] == 1'b1) ? zext_ln1495_fu_324_p1 : data_0_V_read);

assign tmp_289_fu_288_p3 = data_0_V_read[32'd15];

assign tmp_290_fu_302_p3 = data_0_V_read[32'd15];

assign tmp_291_fu_316_p3 = {{xor_ln1495_fu_310_p2}, {10'd0}};

assign tmp_292_fu_342_p3 = data_1_V_read[32'd15];

assign tmp_293_fu_356_p3 = data_1_V_read[32'd15];

assign tmp_294_fu_370_p3 = {{xor_ln1495_95_fu_364_p2}, {10'd0}};

assign tmp_295_fu_396_p3 = data_2_V_read[32'd15];

assign tmp_296_fu_410_p3 = data_2_V_read[32'd15];

assign tmp_297_fu_424_p3 = {{xor_ln1495_96_fu_418_p2}, {10'd0}};

assign tmp_298_fu_450_p3 = data_3_V_read[32'd15];

assign tmp_299_fu_464_p3 = data_3_V_read[32'd15];

assign tmp_300_fu_478_p3 = {{xor_ln1495_97_fu_472_p2}, {10'd0}};

assign tmp_301_fu_504_p3 = data_4_V_read[32'd15];

assign tmp_302_fu_518_p3 = data_4_V_read[32'd15];

assign tmp_303_fu_532_p3 = {{xor_ln1495_98_fu_526_p2}, {10'd0}};

assign tmp_304_fu_558_p3 = data_5_V_read[32'd15];

assign tmp_305_fu_572_p3 = data_5_V_read[32'd15];

assign tmp_306_fu_586_p3 = {{xor_ln1495_99_fu_580_p2}, {10'd0}};

assign tmp_307_fu_612_p3 = data_6_V_read[32'd15];

assign tmp_308_fu_626_p3 = data_6_V_read[32'd15];

assign tmp_309_fu_640_p3 = {{xor_ln1495_100_fu_634_p2}, {10'd0}};

assign tmp_310_fu_666_p3 = data_7_V_read[32'd15];

assign tmp_311_fu_680_p3 = data_7_V_read[32'd15];

assign tmp_312_fu_694_p3 = {{xor_ln1495_101_fu_688_p2}, {10'd0}};

assign tmp_313_fu_720_p3 = data_8_V_read[32'd15];

assign tmp_314_fu_734_p3 = data_8_V_read[32'd15];

assign tmp_315_fu_748_p3 = {{xor_ln1495_102_fu_742_p2}, {10'd0}};

assign tmp_316_fu_774_p3 = data_9_V_read[32'd15];

assign tmp_317_fu_788_p3 = data_9_V_read[32'd15];

assign tmp_318_fu_802_p3 = {{xor_ln1495_103_fu_796_p2}, {10'd0}};

assign tmp_319_fu_828_p3 = data_10_V_read[32'd15];

assign tmp_320_fu_842_p3 = data_10_V_read[32'd15];

assign tmp_321_fu_856_p3 = {{xor_ln1495_104_fu_850_p2}, {10'd0}};

assign tmp_322_fu_882_p3 = data_11_V_read[32'd15];

assign tmp_323_fu_896_p3 = data_11_V_read[32'd15];

assign tmp_324_fu_910_p3 = {{xor_ln1495_105_fu_904_p2}, {10'd0}};

assign tmp_325_fu_936_p3 = data_12_V_read[32'd15];

assign tmp_326_fu_950_p3 = data_12_V_read[32'd15];

assign tmp_327_fu_964_p3 = {{xor_ln1495_106_fu_958_p2}, {10'd0}};

assign tmp_328_fu_990_p3 = data_13_V_read[32'd15];

assign tmp_329_fu_1004_p3 = data_13_V_read[32'd15];

assign tmp_330_fu_1018_p3 = {{xor_ln1495_107_fu_1012_p2}, {10'd0}};

assign tmp_331_fu_1044_p3 = data_14_V_read[32'd15];

assign tmp_332_fu_1058_p3 = data_14_V_read[32'd15];

assign tmp_333_fu_1072_p3 = {{xor_ln1495_108_fu_1066_p2}, {10'd0}};

assign tmp_334_fu_1098_p3 = data_15_V_read[32'd15];

assign tmp_335_fu_1112_p3 = data_15_V_read[32'd15];

assign tmp_336_fu_1126_p3 = {{xor_ln1495_109_fu_1120_p2}, {10'd0}};

assign tmp_337_fu_1152_p3 = data_16_V_read[32'd15];

assign tmp_338_fu_1166_p3 = data_16_V_read[32'd15];

assign tmp_339_fu_1180_p3 = {{xor_ln1495_110_fu_1174_p2}, {10'd0}};

assign tmp_340_fu_1206_p3 = data_17_V_read[32'd15];

assign tmp_341_fu_1220_p3 = data_17_V_read[32'd15];

assign tmp_342_fu_1234_p3 = {{xor_ln1495_111_fu_1228_p2}, {10'd0}};

assign tmp_343_fu_1260_p3 = data_18_V_read[32'd15];

assign tmp_344_fu_1274_p3 = data_18_V_read[32'd15];

assign tmp_345_fu_1288_p3 = {{xor_ln1495_112_fu_1282_p2}, {10'd0}};

assign tmp_346_fu_1314_p3 = data_19_V_read[32'd15];

assign tmp_347_fu_1328_p3 = data_19_V_read[32'd15];

assign tmp_348_fu_1342_p3 = {{xor_ln1495_113_fu_1336_p2}, {10'd0}};

assign tmp_349_fu_1368_p3 = data_20_V_read[32'd15];

assign tmp_350_fu_1382_p3 = data_20_V_read[32'd15];

assign tmp_351_fu_1396_p3 = {{xor_ln1495_114_fu_1390_p2}, {10'd0}};

assign tmp_352_fu_1422_p3 = data_21_V_read[32'd15];

assign tmp_353_fu_1436_p3 = data_21_V_read[32'd15];

assign tmp_354_fu_1450_p3 = {{xor_ln1495_115_fu_1444_p2}, {10'd0}};

assign tmp_355_fu_1476_p3 = data_22_V_read[32'd15];

assign tmp_356_fu_1490_p3 = data_22_V_read[32'd15];

assign tmp_357_fu_1504_p3 = {{xor_ln1495_116_fu_1498_p2}, {10'd0}};

assign tmp_358_fu_1530_p3 = data_23_V_read[32'd15];

assign tmp_359_fu_1544_p3 = data_23_V_read[32'd15];

assign tmp_360_fu_1558_p3 = {{xor_ln1495_117_fu_1552_p2}, {10'd0}};

assign tmp_361_fu_1584_p3 = data_24_V_read[32'd15];

assign tmp_362_fu_1598_p3 = data_24_V_read[32'd15];

assign tmp_363_fu_1612_p3 = {{xor_ln1495_118_fu_1606_p2}, {10'd0}};

assign tmp_364_fu_1638_p3 = data_25_V_read[32'd15];

assign tmp_365_fu_1652_p3 = data_25_V_read[32'd15];

assign tmp_366_fu_1666_p3 = {{xor_ln1495_119_fu_1660_p2}, {10'd0}};

assign tmp_367_fu_1692_p3 = data_26_V_read[32'd15];

assign tmp_368_fu_1706_p3 = data_26_V_read[32'd15];

assign tmp_369_fu_1720_p3 = {{xor_ln1495_120_fu_1714_p2}, {10'd0}};

assign tmp_370_fu_1746_p3 = data_27_V_read[32'd15];

assign tmp_371_fu_1760_p3 = data_27_V_read[32'd15];

assign tmp_372_fu_1774_p3 = {{xor_ln1495_121_fu_1768_p2}, {10'd0}};

assign tmp_373_fu_1800_p3 = data_28_V_read[32'd15];

assign tmp_374_fu_1814_p3 = data_28_V_read[32'd15];

assign tmp_375_fu_1828_p3 = {{xor_ln1495_122_fu_1822_p2}, {10'd0}};

assign tmp_376_fu_1854_p3 = data_29_V_read[32'd15];

assign tmp_377_fu_1868_p3 = data_29_V_read[32'd15];

assign tmp_378_fu_1882_p3 = {{xor_ln1495_123_fu_1876_p2}, {10'd0}};

assign tmp_379_fu_1908_p3 = data_30_V_read[32'd15];

assign tmp_380_fu_1922_p3 = data_30_V_read[32'd15];

assign tmp_381_fu_1936_p3 = {{xor_ln1495_124_fu_1930_p2}, {10'd0}};

assign tmp_382_fu_1962_p3 = data_31_V_read[32'd15];

assign tmp_383_fu_1976_p3 = data_31_V_read[32'd15];

assign tmp_384_fu_1990_p3 = {{xor_ln1495_125_fu_1984_p2}, {10'd0}};

assign xor_ln1495_100_fu_634_p2 = (tmp_308_fu_626_p3 ^ 1'd1);

assign xor_ln1495_101_fu_688_p2 = (tmp_311_fu_680_p3 ^ 1'd1);

assign xor_ln1495_102_fu_742_p2 = (tmp_314_fu_734_p3 ^ 1'd1);

assign xor_ln1495_103_fu_796_p2 = (tmp_317_fu_788_p3 ^ 1'd1);

assign xor_ln1495_104_fu_850_p2 = (tmp_320_fu_842_p3 ^ 1'd1);

assign xor_ln1495_105_fu_904_p2 = (tmp_323_fu_896_p3 ^ 1'd1);

assign xor_ln1495_106_fu_958_p2 = (tmp_326_fu_950_p3 ^ 1'd1);

assign xor_ln1495_107_fu_1012_p2 = (tmp_329_fu_1004_p3 ^ 1'd1);

assign xor_ln1495_108_fu_1066_p2 = (tmp_332_fu_1058_p3 ^ 1'd1);

assign xor_ln1495_109_fu_1120_p2 = (tmp_335_fu_1112_p3 ^ 1'd1);

assign xor_ln1495_110_fu_1174_p2 = (tmp_338_fu_1166_p3 ^ 1'd1);

assign xor_ln1495_111_fu_1228_p2 = (tmp_341_fu_1220_p3 ^ 1'd1);

assign xor_ln1495_112_fu_1282_p2 = (tmp_344_fu_1274_p3 ^ 1'd1);

assign xor_ln1495_113_fu_1336_p2 = (tmp_347_fu_1328_p3 ^ 1'd1);

assign xor_ln1495_114_fu_1390_p2 = (tmp_350_fu_1382_p3 ^ 1'd1);

assign xor_ln1495_115_fu_1444_p2 = (tmp_353_fu_1436_p3 ^ 1'd1);

assign xor_ln1495_116_fu_1498_p2 = (tmp_356_fu_1490_p3 ^ 1'd1);

assign xor_ln1495_117_fu_1552_p2 = (tmp_359_fu_1544_p3 ^ 1'd1);

assign xor_ln1495_118_fu_1606_p2 = (tmp_362_fu_1598_p3 ^ 1'd1);

assign xor_ln1495_119_fu_1660_p2 = (tmp_365_fu_1652_p3 ^ 1'd1);

assign xor_ln1495_120_fu_1714_p2 = (tmp_368_fu_1706_p3 ^ 1'd1);

assign xor_ln1495_121_fu_1768_p2 = (tmp_371_fu_1760_p3 ^ 1'd1);

assign xor_ln1495_122_fu_1822_p2 = (tmp_374_fu_1814_p3 ^ 1'd1);

assign xor_ln1495_123_fu_1876_p2 = (tmp_377_fu_1868_p3 ^ 1'd1);

assign xor_ln1495_124_fu_1930_p2 = (tmp_380_fu_1922_p3 ^ 1'd1);

assign xor_ln1495_125_fu_1984_p2 = (tmp_383_fu_1976_p3 ^ 1'd1);

assign xor_ln1495_95_fu_364_p2 = (tmp_293_fu_356_p3 ^ 1'd1);

assign xor_ln1495_96_fu_418_p2 = (tmp_296_fu_410_p3 ^ 1'd1);

assign xor_ln1495_97_fu_472_p2 = (tmp_299_fu_464_p3 ^ 1'd1);

assign xor_ln1495_98_fu_526_p2 = (tmp_302_fu_518_p3 ^ 1'd1);

assign xor_ln1495_99_fu_580_p2 = (tmp_305_fu_572_p3 ^ 1'd1);

assign xor_ln1495_fu_310_p2 = (tmp_290_fu_302_p3 ^ 1'd1);

assign zext_ln1495_100_fu_648_p1 = tmp_309_fu_640_p3;

assign zext_ln1495_101_fu_702_p1 = tmp_312_fu_694_p3;

assign zext_ln1495_102_fu_756_p1 = tmp_315_fu_748_p3;

assign zext_ln1495_103_fu_810_p1 = tmp_318_fu_802_p3;

assign zext_ln1495_104_fu_864_p1 = tmp_321_fu_856_p3;

assign zext_ln1495_105_fu_918_p1 = tmp_324_fu_910_p3;

assign zext_ln1495_106_fu_972_p1 = tmp_327_fu_964_p3;

assign zext_ln1495_107_fu_1026_p1 = tmp_330_fu_1018_p3;

assign zext_ln1495_108_fu_1080_p1 = tmp_333_fu_1072_p3;

assign zext_ln1495_109_fu_1134_p1 = tmp_336_fu_1126_p3;

assign zext_ln1495_110_fu_1188_p1 = tmp_339_fu_1180_p3;

assign zext_ln1495_111_fu_1242_p1 = tmp_342_fu_1234_p3;

assign zext_ln1495_112_fu_1296_p1 = tmp_345_fu_1288_p3;

assign zext_ln1495_113_fu_1350_p1 = tmp_348_fu_1342_p3;

assign zext_ln1495_114_fu_1404_p1 = tmp_351_fu_1396_p3;

assign zext_ln1495_115_fu_1458_p1 = tmp_354_fu_1450_p3;

assign zext_ln1495_116_fu_1512_p1 = tmp_357_fu_1504_p3;

assign zext_ln1495_117_fu_1566_p1 = tmp_360_fu_1558_p3;

assign zext_ln1495_118_fu_1620_p1 = tmp_363_fu_1612_p3;

assign zext_ln1495_119_fu_1674_p1 = tmp_366_fu_1666_p3;

assign zext_ln1495_120_fu_1728_p1 = tmp_369_fu_1720_p3;

assign zext_ln1495_121_fu_1782_p1 = tmp_372_fu_1774_p3;

assign zext_ln1495_122_fu_1836_p1 = tmp_375_fu_1828_p3;

assign zext_ln1495_123_fu_1890_p1 = tmp_378_fu_1882_p3;

assign zext_ln1495_124_fu_1944_p1 = tmp_381_fu_1936_p3;

assign zext_ln1495_125_fu_1998_p1 = tmp_384_fu_1990_p3;

assign zext_ln1495_95_fu_378_p1 = tmp_294_fu_370_p3;

assign zext_ln1495_96_fu_432_p1 = tmp_297_fu_424_p3;

assign zext_ln1495_97_fu_486_p1 = tmp_300_fu_478_p3;

assign zext_ln1495_98_fu_540_p1 = tmp_303_fu_532_p3;

assign zext_ln1495_99_fu_594_p1 = tmp_306_fu_586_p3;

assign zext_ln1495_fu_324_p1 = tmp_291_fu_316_p3;

endmodule //relu_max_ap_fixed_ap_fixed_1_relu1_config13_s
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module relu_max_ap_fixed_ap_fixed_1_relu1_config5_s (
        ap_ready,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        data_32_V_read,
        data_33_V_read,
        data_34_V_read,
        data_35_V_read,
        data_36_V_read,
        data_37_V_read,
        data_38_V_read,
        data_39_V_read,
        data_40_V_read,
        data_41_V_read,
        data_42_V_read,
        data_43_V_read,
        data_44_V_read,
        data_45_V_read,
        data_46_V_read,
        data_47_V_read,
        data_48_V_read,
        data_49_V_read,
        data_50_V_read,
        data_51_V_read,
        data_52_V_read,
        data_53_V_read,
        data_54_V_read,
        data_55_V_read,
        data_56_V_read,
        data_57_V_read,
        data_58_V_read,
        data_59_V_read,
        data_60_V_read,
        data_61_V_read,
        data_62_V_read,
        data_63_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63
);


output   ap_ready;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
input  [15:0] data_32_V_read;
input  [15:0] data_33_V_read;
input  [15:0] data_34_V_read;
input  [15:0] data_35_V_read;
input  [15:0] data_36_V_read;
input  [15:0] data_37_V_read;
input  [15:0] data_38_V_read;
input  [15:0] data_39_V_read;
input  [15:0] data_40_V_read;
input  [15:0] data_41_V_read;
input  [15:0] data_42_V_read;
input  [15:0] data_43_V_read;
input  [15:0] data_44_V_read;
input  [15:0] data_45_V_read;
input  [15:0] data_46_V_read;
input  [15:0] data_47_V_read;
input  [15:0] data_48_V_read;
input  [15:0] data_49_V_read;
input  [15:0] data_50_V_read;
input  [15:0] data_51_V_read;
input  [15:0] data_52_V_read;
input  [15:0] data_53_V_read;
input  [15:0] data_54_V_read;
input  [15:0] data_55_V_read;
input  [15:0] data_56_V_read;
input  [15:0] data_57_V_read;
input  [15:0] data_58_V_read;
input  [15:0] data_59_V_read;
input  [15:0] data_60_V_read;
input  [15:0] data_61_V_read;
input  [15:0] data_62_V_read;
input  [15:0] data_63_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
output  [15:0] ap_return_32;
output  [15:0] ap_return_33;
output  [15:0] ap_return_34;
output  [15:0] ap_return_35;
output  [15:0] ap_return_36;
output  [15:0] ap_return_37;
output  [15:0] ap_return_38;
output  [15:0] ap_return_39;
output  [15:0] ap_return_40;
output  [15:0] ap_return_41;
output  [15:0] ap_return_42;
output  [15:0] ap_return_43;
output  [15:0] ap_return_44;
output  [15:0] ap_return_45;
output  [15:0] ap_return_46;
output  [15:0] ap_return_47;
output  [15:0] ap_return_48;
output  [15:0] ap_return_49;
output  [15:0] ap_return_50;
output  [15:0] ap_return_51;
output  [15:0] ap_return_52;
output  [15:0] ap_return_53;
output  [15:0] ap_return_54;
output  [15:0] ap_return_55;
output  [15:0] ap_return_56;
output  [15:0] ap_return_57;
output  [15:0] ap_return_58;
output  [15:0] ap_return_59;
output  [15:0] ap_return_60;
output  [15:0] ap_return_61;
output  [15:0] ap_return_62;
output  [15:0] ap_return_63;

wire   [0:0] tmp_98_fu_558_p3;
wire   [0:0] xor_ln1495_fu_566_p2;
wire   [10:0] tmp_99_fu_572_p3;
wire   [0:0] tmp_97_fu_544_p3;
wire   [0:0] icmp_ln1494_fu_552_p2;
wire   [0:0] or_ln1495_fu_584_p2;
wire   [15:0] zext_ln1495_fu_580_p1;
wire   [0:0] tmp_101_fu_612_p3;
wire   [0:0] xor_ln1495_32_fu_620_p2;
wire   [10:0] tmp_102_fu_626_p3;
wire   [0:0] tmp_100_fu_598_p3;
wire   [0:0] icmp_ln1494_1_fu_606_p2;
wire   [0:0] or_ln1495_32_fu_638_p2;
wire   [15:0] zext_ln1495_32_fu_634_p1;
wire   [0:0] tmp_104_fu_666_p3;
wire   [0:0] xor_ln1495_33_fu_674_p2;
wire   [10:0] tmp_105_fu_680_p3;
wire   [0:0] tmp_103_fu_652_p3;
wire   [0:0] icmp_ln1494_2_fu_660_p2;
wire   [0:0] or_ln1495_33_fu_692_p2;
wire   [15:0] zext_ln1495_33_fu_688_p1;
wire   [0:0] tmp_107_fu_720_p3;
wire   [0:0] xor_ln1495_34_fu_728_p2;
wire   [10:0] tmp_108_fu_734_p3;
wire   [0:0] tmp_106_fu_706_p3;
wire   [0:0] icmp_ln1494_3_fu_714_p2;
wire   [0:0] or_ln1495_34_fu_746_p2;
wire   [15:0] zext_ln1495_34_fu_742_p1;
wire   [0:0] tmp_110_fu_774_p3;
wire   [0:0] xor_ln1495_35_fu_782_p2;
wire   [10:0] tmp_111_fu_788_p3;
wire   [0:0] tmp_109_fu_760_p3;
wire   [0:0] icmp_ln1494_4_fu_768_p2;
wire   [0:0] or_ln1495_35_fu_800_p2;
wire   [15:0] zext_ln1495_35_fu_796_p1;
wire   [0:0] tmp_113_fu_828_p3;
wire   [0:0] xor_ln1495_36_fu_836_p2;
wire   [10:0] tmp_114_fu_842_p3;
wire   [0:0] tmp_112_fu_814_p3;
wire   [0:0] icmp_ln1494_5_fu_822_p2;
wire   [0:0] or_ln1495_36_fu_854_p2;
wire   [15:0] zext_ln1495_36_fu_850_p1;
wire   [0:0] tmp_116_fu_882_p3;
wire   [0:0] xor_ln1495_37_fu_890_p2;
wire   [10:0] tmp_117_fu_896_p3;
wire   [0:0] tmp_115_fu_868_p3;
wire   [0:0] icmp_ln1494_6_fu_876_p2;
wire   [0:0] or_ln1495_37_fu_908_p2;
wire   [15:0] zext_ln1495_37_fu_904_p1;
wire   [0:0] tmp_119_fu_936_p3;
wire   [0:0] xor_ln1495_38_fu_944_p2;
wire   [10:0] tmp_120_fu_950_p3;
wire   [0:0] tmp_118_fu_922_p3;
wire   [0:0] icmp_ln1494_7_fu_930_p2;
wire   [0:0] or_ln1495_38_fu_962_p2;
wire   [15:0] zext_ln1495_38_fu_958_p1;
wire   [0:0] tmp_122_fu_990_p3;
wire   [0:0] xor_ln1495_39_fu_998_p2;
wire   [10:0] tmp_123_fu_1004_p3;
wire   [0:0] tmp_121_fu_976_p3;
wire   [0:0] icmp_ln1494_8_fu_984_p2;
wire   [0:0] or_ln1495_39_fu_1016_p2;
wire   [15:0] zext_ln1495_39_fu_1012_p1;
wire   [0:0] tmp_125_fu_1044_p3;
wire   [0:0] xor_ln1495_40_fu_1052_p2;
wire   [10:0] tmp_126_fu_1058_p3;
wire   [0:0] tmp_124_fu_1030_p3;
wire   [0:0] icmp_ln1494_9_fu_1038_p2;
wire   [0:0] or_ln1495_40_fu_1070_p2;
wire   [15:0] zext_ln1495_40_fu_1066_p1;
wire   [0:0] tmp_128_fu_1098_p3;
wire   [0:0] xor_ln1495_41_fu_1106_p2;
wire   [10:0] tmp_129_fu_1112_p3;
wire   [0:0] tmp_127_fu_1084_p3;
wire   [0:0] icmp_ln1494_10_fu_1092_p2;
wire   [0:0] or_ln1495_41_fu_1124_p2;
wire   [15:0] zext_ln1495_41_fu_1120_p1;
wire   [0:0] tmp_131_fu_1152_p3;
wire   [0:0] xor_ln1495_42_fu_1160_p2;
wire   [10:0] tmp_132_fu_1166_p3;
wire   [0:0] tmp_130_fu_1138_p3;
wire   [0:0] icmp_ln1494_11_fu_1146_p2;
wire   [0:0] or_ln1495_42_fu_1178_p2;
wire   [15:0] zext_ln1495_42_fu_1174_p1;
wire   [0:0] tmp_134_fu_1206_p3;
wire   [0:0] xor_ln1495_43_fu_1214_p2;
wire   [10:0] tmp_135_fu_1220_p3;
wire   [0:0] tmp_133_fu_1192_p3;
wire   [0:0] icmp_ln1494_12_fu_1200_p2;
wire   [0:0] or_ln1495_43_fu_1232_p2;
wire   [15:0] zext_ln1495_43_fu_1228_p1;
wire   [0:0] tmp_137_fu_1260_p3;
wire   [0:0] xor_ln1495_44_fu_1268_p2;
wire   [10:0] tmp_138_fu_1274_p3;
wire   [0:0] tmp_136_fu_1246_p3;
wire   [0:0] icmp_ln1494_13_fu_1254_p2;
wire   [0:0] or_ln1495_44_fu_1286_p2;
wire   [15:0] zext_ln1495_44_fu_1282_p1;
wire   [0:0] tmp_140_fu_1314_p3;
wire   [0:0] xor_ln1495_45_fu_1322_p2;
wire   [10:0] tmp_141_fu_1328_p3;
wire   [0:0] tmp_139_fu_1300_p3;
wire   [0:0] icmp_ln1494_14_fu_1308_p2;
wire   [0:0] or_ln1495_45_fu_1340_p2;
wire   [15:0] zext_ln1495_45_fu_1336_p1;
wire   [0:0] tmp_143_fu_1368_p3;
wire   [0:0] xor_ln1495_46_fu_1376_p2;
wire   [10:0] tmp_144_fu_1382_p3;
wire   [0:0] tmp_142_fu_1354_p3;
wire   [0:0] icmp_ln1494_15_fu_1362_p2;
wire   [0:0] or_ln1495_46_fu_1394_p2;
wire   [15:0] zext_ln1495_46_fu_1390_p1;
wire   [0:0] tmp_146_fu_1422_p3;
wire   [0:0] xor_ln1495_47_fu_1430_p2;
wire   [10:0] tmp_147_fu_1436_p3;
wire   [0:0] tmp_145_fu_1408_p3;
wire   [0:0] icmp_ln1494_16_fu_1416_p2;
wire   [0:0] or_ln1495_47_fu_1448_p2;
wire   [15:0] zext_ln1495_47_fu_1444_p1;
wire   [0:0] tmp_149_fu_1476_p3;
wire   [0:0] xor_ln1495_48_fu_1484_p2;
wire   [10:0] tmp_150_fu_1490_p3;
wire   [0:0] tmp_148_fu_1462_p3;
wire   [0:0] icmp_ln1494_17_fu_1470_p2;
wire   [0:0] or_ln1495_48_fu_1502_p2;
wire   [15:0] zext_ln1495_48_fu_1498_p1;
wire   [0:0] tmp_152_fu_1530_p3;
wire   [0:0] xor_ln1495_49_fu_1538_p2;
wire   [10:0] tmp_153_fu_1544_p3;
wire   [0:0] tmp_151_fu_1516_p3;
wire   [0:0] icmp_ln1494_18_fu_1524_p2;
wire   [0:0] or_ln1495_49_fu_1556_p2;
wire   [15:0] zext_ln1495_49_fu_1552_p1;
wire   [0:0] tmp_155_fu_1584_p3;
wire   [0:0] xor_ln1495_50_fu_1592_p2;
wire   [10:0] tmp_156_fu_1598_p3;
wire   [0:0] tmp_154_fu_1570_p3;
wire   [0:0] icmp_ln1494_19_fu_1578_p2;
wire   [0:0] or_ln1495_50_fu_1610_p2;
wire   [15:0] zext_ln1495_50_fu_1606_p1;
wire   [0:0] tmp_158_fu_1638_p3;
wire   [0:0] xor_ln1495_51_fu_1646_p2;
wire   [10:0] tmp_159_fu_1652_p3;
wire   [0:0] tmp_157_fu_1624_p3;
wire   [0:0] icmp_ln1494_20_fu_1632_p2;
wire   [0:0] or_ln1495_51_fu_1664_p2;
wire   [15:0] zext_ln1495_51_fu_1660_p1;
wire   [0:0] tmp_161_fu_1692_p3;
wire   [0:0] xor_ln1495_52_fu_1700_p2;
wire   [10:0] tmp_162_fu_1706_p3;
wire   [0:0] tmp_160_fu_1678_p3;
wire   [0:0] icmp_ln1494_21_fu_1686_p2;
wire   [0:0] or_ln1495_52_fu_1718_p2;
wire   [15:0] zext_ln1495_52_fu_1714_p1;
wire   [0:0] tmp_164_fu_1746_p3;
wire   [0:0] xor_ln1495_53_fu_1754_p2;
wire   [10:0] tmp_165_fu_1760_p3;
wire   [0:0] tmp_163_fu_1732_p3;
wire   [0:0] icmp_ln1494_22_fu_1740_p2;
wire   [0:0] or_ln1495_53_fu_1772_p2;
wire   [15:0] zext_ln1495_53_fu_1768_p1;
wire   [0:0] tmp_167_fu_1800_p3;
wire   [0:0] xor_ln1495_54_fu_1808_p2;
wire   [10:0] tmp_168_fu_1814_p3;
wire   [0:0] tmp_166_fu_1786_p3;
wire   [0:0] icmp_ln1494_23_fu_1794_p2;
wire   [0:0] or_ln1495_54_fu_1826_p2;
wire   [15:0] zext_ln1495_54_fu_1822_p1;
wire   [0:0] tmp_170_fu_1854_p3;
wire   [0:0] xor_ln1495_55_fu_1862_p2;
wire   [10:0] tmp_171_fu_1868_p3;
wire   [0:0] tmp_169_fu_1840_p3;
wire   [0:0] icmp_ln1494_24_fu_1848_p2;
wire   [0:0] or_ln1495_55_fu_1880_p2;
wire   [15:0] zext_ln1495_55_fu_1876_p1;
wire   [0:0] tmp_173_fu_1908_p3;
wire   [0:0] xor_ln1495_56_fu_1916_p2;
wire   [10:0] tmp_174_fu_1922_p3;
wire   [0:0] tmp_172_fu_1894_p3;
wire   [0:0] icmp_ln1494_25_fu_1902_p2;
wire   [0:0] or_ln1495_56_fu_1934_p2;
wire   [15:0] zext_ln1495_56_fu_1930_p1;
wire   [0:0] tmp_176_fu_1962_p3;
wire   [0:0] xor_ln1495_57_fu_1970_p2;
wire   [10:0] tmp_177_fu_1976_p3;
wire   [0:0] tmp_175_fu_1948_p3;
wire   [0:0] icmp_ln1494_26_fu_1956_p2;
wire   [0:0] or_ln1495_57_fu_1988_p2;
wire   [15:0] zext_ln1495_57_fu_1984_p1;
wire   [0:0] tmp_179_fu_2016_p3;
wire   [0:0] xor_ln1495_58_fu_2024_p2;
wire   [10:0] tmp_180_fu_2030_p3;
wire   [0:0] tmp_178_fu_2002_p3;
wire   [0:0] icmp_ln1494_27_fu_2010_p2;
wire   [0:0] or_ln1495_58_fu_2042_p2;
wire   [15:0] zext_ln1495_58_fu_2038_p1;
wire   [0:0] tmp_182_fu_2070_p3;
wire   [0:0] xor_ln1495_59_fu_2078_p2;
wire   [10:0] tmp_183_fu_2084_p3;
wire   [0:0] tmp_181_fu_2056_p3;
wire   [0:0] icmp_ln1494_28_fu_2064_p2;
wire   [0:0] or_ln1495_59_fu_2096_p2;
wire   [15:0] zext_ln1495_59_fu_2092_p1;
wire   [0:0] tmp_185_fu_2124_p3;
wire   [0:0] xor_ln1495_60_fu_2132_p2;
wire   [10:0] tmp_186_fu_2138_p3;
wire   [0:0] tmp_184_fu_2110_p3;
wire   [0:0] icmp_ln1494_29_fu_2118_p2;
wire   [0:0] or_ln1495_60_fu_2150_p2;
wire   [15:0] zext_ln1495_60_fu_2146_p1;
wire   [0:0] tmp_188_fu_2178_p3;
wire   [0:0] xor_ln1495_61_fu_2186_p2;
wire   [10:0] tmp_189_fu_2192_p3;
wire   [0:0] tmp_187_fu_2164_p3;
wire   [0:0] icmp_ln1494_30_fu_2172_p2;
wire   [0:0] or_ln1495_61_fu_2204_p2;
wire   [15:0] zext_ln1495_61_fu_2200_p1;
wire   [0:0] tmp_191_fu_2232_p3;
wire   [0:0] xor_ln1495_62_fu_2240_p2;
wire   [10:0] tmp_192_fu_2246_p3;
wire   [0:0] tmp_190_fu_2218_p3;
wire   [0:0] icmp_ln1494_31_fu_2226_p2;
wire   [0:0] or_ln1495_62_fu_2258_p2;
wire   [15:0] zext_ln1495_62_fu_2254_p1;
wire   [0:0] tmp_194_fu_2286_p3;
wire   [0:0] xor_ln1495_63_fu_2294_p2;
wire   [10:0] tmp_195_fu_2300_p3;
wire   [0:0] tmp_193_fu_2272_p3;
wire   [0:0] icmp_ln1494_32_fu_2280_p2;
wire   [0:0] or_ln1495_63_fu_2312_p2;
wire   [15:0] zext_ln1495_63_fu_2308_p1;
wire   [0:0] tmp_197_fu_2340_p3;
wire   [0:0] xor_ln1495_64_fu_2348_p2;
wire   [10:0] tmp_198_fu_2354_p3;
wire   [0:0] tmp_196_fu_2326_p3;
wire   [0:0] icmp_ln1494_33_fu_2334_p2;
wire   [0:0] or_ln1495_64_fu_2366_p2;
wire   [15:0] zext_ln1495_64_fu_2362_p1;
wire   [0:0] tmp_200_fu_2394_p3;
wire   [0:0] xor_ln1495_65_fu_2402_p2;
wire   [10:0] tmp_201_fu_2408_p3;
wire   [0:0] tmp_199_fu_2380_p3;
wire   [0:0] icmp_ln1494_34_fu_2388_p2;
wire   [0:0] or_ln1495_65_fu_2420_p2;
wire   [15:0] zext_ln1495_65_fu_2416_p1;
wire   [0:0] tmp_203_fu_2448_p3;
wire   [0:0] xor_ln1495_66_fu_2456_p2;
wire   [10:0] tmp_204_fu_2462_p3;
wire   [0:0] tmp_202_fu_2434_p3;
wire   [0:0] icmp_ln1494_35_fu_2442_p2;
wire   [0:0] or_ln1495_66_fu_2474_p2;
wire   [15:0] zext_ln1495_66_fu_2470_p1;
wire   [0:0] tmp_206_fu_2502_p3;
wire   [0:0] xor_ln1495_67_fu_2510_p2;
wire   [10:0] tmp_207_fu_2516_p3;
wire   [0:0] tmp_205_fu_2488_p3;
wire   [0:0] icmp_ln1494_36_fu_2496_p2;
wire   [0:0] or_ln1495_67_fu_2528_p2;
wire   [15:0] zext_ln1495_67_fu_2524_p1;
wire   [0:0] tmp_209_fu_2556_p3;
wire   [0:0] xor_ln1495_68_fu_2564_p2;
wire   [10:0] tmp_210_fu_2570_p3;
wire   [0:0] tmp_208_fu_2542_p3;
wire   [0:0] icmp_ln1494_37_fu_2550_p2;
wire   [0:0] or_ln1495_68_fu_2582_p2;
wire   [15:0] zext_ln1495_68_fu_2578_p1;
wire   [0:0] tmp_212_fu_2610_p3;
wire   [0:0] xor_ln1495_69_fu_2618_p2;
wire   [10:0] tmp_213_fu_2624_p3;
wire   [0:0] tmp_211_fu_2596_p3;
wire   [0:0] icmp_ln1494_38_fu_2604_p2;
wire   [0:0] or_ln1495_69_fu_2636_p2;
wire   [15:0] zext_ln1495_69_fu_2632_p1;
wire   [0:0] tmp_215_fu_2664_p3;
wire   [0:0] xor_ln1495_70_fu_2672_p2;
wire   [10:0] tmp_216_fu_2678_p3;
wire   [0:0] tmp_214_fu_2650_p3;
wire   [0:0] icmp_ln1494_39_fu_2658_p2;
wire   [0:0] or_ln1495_70_fu_2690_p2;
wire   [15:0] zext_ln1495_70_fu_2686_p1;
wire   [0:0] tmp_218_fu_2718_p3;
wire   [0:0] xor_ln1495_71_fu_2726_p2;
wire   [10:0] tmp_219_fu_2732_p3;
wire   [0:0] tmp_217_fu_2704_p3;
wire   [0:0] icmp_ln1494_40_fu_2712_p2;
wire   [0:0] or_ln1495_71_fu_2744_p2;
wire   [15:0] zext_ln1495_71_fu_2740_p1;
wire   [0:0] tmp_221_fu_2772_p3;
wire   [0:0] xor_ln1495_72_fu_2780_p2;
wire   [10:0] tmp_222_fu_2786_p3;
wire   [0:0] tmp_220_fu_2758_p3;
wire   [0:0] icmp_ln1494_41_fu_2766_p2;
wire   [0:0] or_ln1495_72_fu_2798_p2;
wire   [15:0] zext_ln1495_72_fu_2794_p1;
wire   [0:0] tmp_224_fu_2826_p3;
wire   [0:0] xor_ln1495_73_fu_2834_p2;
wire   [10:0] tmp_225_fu_2840_p3;
wire   [0:0] tmp_223_fu_2812_p3;
wire   [0:0] icmp_ln1494_42_fu_2820_p2;
wire   [0:0] or_ln1495_73_fu_2852_p2;
wire   [15:0] zext_ln1495_73_fu_2848_p1;
wire   [0:0] tmp_227_fu_2880_p3;
wire   [0:0] xor_ln1495_74_fu_2888_p2;
wire   [10:0] tmp_228_fu_2894_p3;
wire   [0:0] tmp_226_fu_2866_p3;
wire   [0:0] icmp_ln1494_43_fu_2874_p2;
wire   [0:0] or_ln1495_74_fu_2906_p2;
wire   [15:0] zext_ln1495_74_fu_2902_p1;
wire   [0:0] tmp_230_fu_2934_p3;
wire   [0:0] xor_ln1495_75_fu_2942_p2;
wire   [10:0] tmp_231_fu_2948_p3;
wire   [0:0] tmp_229_fu_2920_p3;
wire   [0:0] icmp_ln1494_44_fu_2928_p2;
wire   [0:0] or_ln1495_75_fu_2960_p2;
wire   [15:0] zext_ln1495_75_fu_2956_p1;
wire   [0:0] tmp_233_fu_2988_p3;
wire   [0:0] xor_ln1495_76_fu_2996_p2;
wire   [10:0] tmp_234_fu_3002_p3;
wire   [0:0] tmp_232_fu_2974_p3;
wire   [0:0] icmp_ln1494_45_fu_2982_p2;
wire   [0:0] or_ln1495_76_fu_3014_p2;
wire   [15:0] zext_ln1495_76_fu_3010_p1;
wire   [0:0] tmp_236_fu_3042_p3;
wire   [0:0] xor_ln1495_77_fu_3050_p2;
wire   [10:0] tmp_237_fu_3056_p3;
wire   [0:0] tmp_235_fu_3028_p3;
wire   [0:0] icmp_ln1494_46_fu_3036_p2;
wire   [0:0] or_ln1495_77_fu_3068_p2;
wire   [15:0] zext_ln1495_77_fu_3064_p1;
wire   [0:0] tmp_239_fu_3096_p3;
wire   [0:0] xor_ln1495_78_fu_3104_p2;
wire   [10:0] tmp_240_fu_3110_p3;
wire   [0:0] tmp_238_fu_3082_p3;
wire   [0:0] icmp_ln1494_47_fu_3090_p2;
wire   [0:0] or_ln1495_78_fu_3122_p2;
wire   [15:0] zext_ln1495_78_fu_3118_p1;
wire   [0:0] tmp_242_fu_3150_p3;
wire   [0:0] xor_ln1495_79_fu_3158_p2;
wire   [10:0] tmp_243_fu_3164_p3;
wire   [0:0] tmp_241_fu_3136_p3;
wire   [0:0] icmp_ln1494_48_fu_3144_p2;
wire   [0:0] or_ln1495_79_fu_3176_p2;
wire   [15:0] zext_ln1495_79_fu_3172_p1;
wire   [0:0] tmp_245_fu_3204_p3;
wire   [0:0] xor_ln1495_80_fu_3212_p2;
wire   [10:0] tmp_246_fu_3218_p3;
wire   [0:0] tmp_244_fu_3190_p3;
wire   [0:0] icmp_ln1494_49_fu_3198_p2;
wire   [0:0] or_ln1495_80_fu_3230_p2;
wire   [15:0] zext_ln1495_80_fu_3226_p1;
wire   [0:0] tmp_248_fu_3258_p3;
wire   [0:0] xor_ln1495_81_fu_3266_p2;
wire   [10:0] tmp_249_fu_3272_p3;
wire   [0:0] tmp_247_fu_3244_p3;
wire   [0:0] icmp_ln1494_50_fu_3252_p2;
wire   [0:0] or_ln1495_81_fu_3284_p2;
wire   [15:0] zext_ln1495_81_fu_3280_p1;
wire   [0:0] tmp_251_fu_3312_p3;
wire   [0:0] xor_ln1495_82_fu_3320_p2;
wire   [10:0] tmp_252_fu_3326_p3;
wire   [0:0] tmp_250_fu_3298_p3;
wire   [0:0] icmp_ln1494_51_fu_3306_p2;
wire   [0:0] or_ln1495_82_fu_3338_p2;
wire   [15:0] zext_ln1495_82_fu_3334_p1;
wire   [0:0] tmp_254_fu_3366_p3;
wire   [0:0] xor_ln1495_83_fu_3374_p2;
wire   [10:0] tmp_255_fu_3380_p3;
wire   [0:0] tmp_253_fu_3352_p3;
wire   [0:0] icmp_ln1494_52_fu_3360_p2;
wire   [0:0] or_ln1495_83_fu_3392_p2;
wire   [15:0] zext_ln1495_83_fu_3388_p1;
wire   [0:0] tmp_257_fu_3420_p3;
wire   [0:0] xor_ln1495_84_fu_3428_p2;
wire   [10:0] tmp_258_fu_3434_p3;
wire   [0:0] tmp_256_fu_3406_p3;
wire   [0:0] icmp_ln1494_53_fu_3414_p2;
wire   [0:0] or_ln1495_84_fu_3446_p2;
wire   [15:0] zext_ln1495_84_fu_3442_p1;
wire   [0:0] tmp_260_fu_3474_p3;
wire   [0:0] xor_ln1495_85_fu_3482_p2;
wire   [10:0] tmp_261_fu_3488_p3;
wire   [0:0] tmp_259_fu_3460_p3;
wire   [0:0] icmp_ln1494_54_fu_3468_p2;
wire   [0:0] or_ln1495_85_fu_3500_p2;
wire   [15:0] zext_ln1495_85_fu_3496_p1;
wire   [0:0] tmp_263_fu_3528_p3;
wire   [0:0] xor_ln1495_86_fu_3536_p2;
wire   [10:0] tmp_264_fu_3542_p3;
wire   [0:0] tmp_262_fu_3514_p3;
wire   [0:0] icmp_ln1494_55_fu_3522_p2;
wire   [0:0] or_ln1495_86_fu_3554_p2;
wire   [15:0] zext_ln1495_86_fu_3550_p1;
wire   [0:0] tmp_266_fu_3582_p3;
wire   [0:0] xor_ln1495_87_fu_3590_p2;
wire   [10:0] tmp_267_fu_3596_p3;
wire   [0:0] tmp_265_fu_3568_p3;
wire   [0:0] icmp_ln1494_56_fu_3576_p2;
wire   [0:0] or_ln1495_87_fu_3608_p2;
wire   [15:0] zext_ln1495_87_fu_3604_p1;
wire   [0:0] tmp_269_fu_3636_p3;
wire   [0:0] xor_ln1495_88_fu_3644_p2;
wire   [10:0] tmp_270_fu_3650_p3;
wire   [0:0] tmp_268_fu_3622_p3;
wire   [0:0] icmp_ln1494_57_fu_3630_p2;
wire   [0:0] or_ln1495_88_fu_3662_p2;
wire   [15:0] zext_ln1495_88_fu_3658_p1;
wire   [0:0] tmp_272_fu_3690_p3;
wire   [0:0] xor_ln1495_89_fu_3698_p2;
wire   [10:0] tmp_273_fu_3704_p3;
wire   [0:0] tmp_271_fu_3676_p3;
wire   [0:0] icmp_ln1494_58_fu_3684_p2;
wire   [0:0] or_ln1495_89_fu_3716_p2;
wire   [15:0] zext_ln1495_89_fu_3712_p1;
wire   [0:0] tmp_275_fu_3744_p3;
wire   [0:0] xor_ln1495_90_fu_3752_p2;
wire   [10:0] tmp_276_fu_3758_p3;
wire   [0:0] tmp_274_fu_3730_p3;
wire   [0:0] icmp_ln1494_59_fu_3738_p2;
wire   [0:0] or_ln1495_90_fu_3770_p2;
wire   [15:0] zext_ln1495_90_fu_3766_p1;
wire   [0:0] tmp_278_fu_3798_p3;
wire   [0:0] xor_ln1495_91_fu_3806_p2;
wire   [10:0] tmp_279_fu_3812_p3;
wire   [0:0] tmp_277_fu_3784_p3;
wire   [0:0] icmp_ln1494_60_fu_3792_p2;
wire   [0:0] or_ln1495_91_fu_3824_p2;
wire   [15:0] zext_ln1495_91_fu_3820_p1;
wire   [0:0] tmp_281_fu_3852_p3;
wire   [0:0] xor_ln1495_92_fu_3860_p2;
wire   [10:0] tmp_282_fu_3866_p3;
wire   [0:0] tmp_280_fu_3838_p3;
wire   [0:0] icmp_ln1494_61_fu_3846_p2;
wire   [0:0] or_ln1495_92_fu_3878_p2;
wire   [15:0] zext_ln1495_92_fu_3874_p1;
wire   [0:0] tmp_284_fu_3906_p3;
wire   [0:0] xor_ln1495_93_fu_3914_p2;
wire   [10:0] tmp_285_fu_3920_p3;
wire   [0:0] tmp_283_fu_3892_p3;
wire   [0:0] icmp_ln1494_62_fu_3900_p2;
wire   [0:0] or_ln1495_93_fu_3932_p2;
wire   [15:0] zext_ln1495_93_fu_3928_p1;
wire   [0:0] tmp_287_fu_3960_p3;
wire   [0:0] xor_ln1495_94_fu_3968_p2;
wire   [10:0] tmp_288_fu_3974_p3;
wire   [0:0] tmp_286_fu_3946_p3;
wire   [0:0] icmp_ln1494_63_fu_3954_p2;
wire   [0:0] or_ln1495_94_fu_3986_p2;
wire   [15:0] zext_ln1495_94_fu_3982_p1;
wire   [15:0] select_ln1495_fu_590_p3;
wire   [15:0] select_ln1495_32_fu_644_p3;
wire   [15:0] select_ln1495_33_fu_698_p3;
wire   [15:0] select_ln1495_34_fu_752_p3;
wire   [15:0] select_ln1495_35_fu_806_p3;
wire   [15:0] select_ln1495_36_fu_860_p3;
wire   [15:0] select_ln1495_37_fu_914_p3;
wire   [15:0] select_ln1495_38_fu_968_p3;
wire   [15:0] select_ln1495_39_fu_1022_p3;
wire   [15:0] select_ln1495_40_fu_1076_p3;
wire   [15:0] select_ln1495_41_fu_1130_p3;
wire   [15:0] select_ln1495_42_fu_1184_p3;
wire   [15:0] select_ln1495_43_fu_1238_p3;
wire   [15:0] select_ln1495_44_fu_1292_p3;
wire   [15:0] select_ln1495_45_fu_1346_p3;
wire   [15:0] select_ln1495_46_fu_1400_p3;
wire   [15:0] select_ln1495_47_fu_1454_p3;
wire   [15:0] select_ln1495_48_fu_1508_p3;
wire   [15:0] select_ln1495_49_fu_1562_p3;
wire   [15:0] select_ln1495_50_fu_1616_p3;
wire   [15:0] select_ln1495_51_fu_1670_p3;
wire   [15:0] select_ln1495_52_fu_1724_p3;
wire   [15:0] select_ln1495_53_fu_1778_p3;
wire   [15:0] select_ln1495_54_fu_1832_p3;
wire   [15:0] select_ln1495_55_fu_1886_p3;
wire   [15:0] select_ln1495_56_fu_1940_p3;
wire   [15:0] select_ln1495_57_fu_1994_p3;
wire   [15:0] select_ln1495_58_fu_2048_p3;
wire   [15:0] select_ln1495_59_fu_2102_p3;
wire   [15:0] select_ln1495_60_fu_2156_p3;
wire   [15:0] select_ln1495_61_fu_2210_p3;
wire   [15:0] select_ln1495_62_fu_2264_p3;
wire   [15:0] select_ln1495_63_fu_2318_p3;
wire   [15:0] select_ln1495_64_fu_2372_p3;
wire   [15:0] select_ln1495_65_fu_2426_p3;
wire   [15:0] select_ln1495_66_fu_2480_p3;
wire   [15:0] select_ln1495_67_fu_2534_p3;
wire   [15:0] select_ln1495_68_fu_2588_p3;
wire   [15:0] select_ln1495_69_fu_2642_p3;
wire   [15:0] select_ln1495_70_fu_2696_p3;
wire   [15:0] select_ln1495_71_fu_2750_p3;
wire   [15:0] select_ln1495_72_fu_2804_p3;
wire   [15:0] select_ln1495_73_fu_2858_p3;
wire   [15:0] select_ln1495_74_fu_2912_p3;
wire   [15:0] select_ln1495_75_fu_2966_p3;
wire   [15:0] select_ln1495_76_fu_3020_p3;
wire   [15:0] select_ln1495_77_fu_3074_p3;
wire   [15:0] select_ln1495_78_fu_3128_p3;
wire   [15:0] select_ln1495_79_fu_3182_p3;
wire   [15:0] select_ln1495_80_fu_3236_p3;
wire   [15:0] select_ln1495_81_fu_3290_p3;
wire   [15:0] select_ln1495_82_fu_3344_p3;
wire   [15:0] select_ln1495_83_fu_3398_p3;
wire   [15:0] select_ln1495_84_fu_3452_p3;
wire   [15:0] select_ln1495_85_fu_3506_p3;
wire   [15:0] select_ln1495_86_fu_3560_p3;
wire   [15:0] select_ln1495_87_fu_3614_p3;
wire   [15:0] select_ln1495_88_fu_3668_p3;
wire   [15:0] select_ln1495_89_fu_3722_p3;
wire   [15:0] select_ln1495_90_fu_3776_p3;
wire   [15:0] select_ln1495_91_fu_3830_p3;
wire   [15:0] select_ln1495_92_fu_3884_p3;
wire   [15:0] select_ln1495_93_fu_3938_p3;
wire   [15:0] select_ln1495_94_fu_3992_p3;

assign ap_ready = 1'b1;

assign ap_return_0 = select_ln1495_fu_590_p3;

assign ap_return_1 = select_ln1495_32_fu_644_p3;

assign ap_return_10 = select_ln1495_41_fu_1130_p3;

assign ap_return_11 = select_ln1495_42_fu_1184_p3;

assign ap_return_12 = select_ln1495_43_fu_1238_p3;

assign ap_return_13 = select_ln1495_44_fu_1292_p3;

assign ap_return_14 = select_ln1495_45_fu_1346_p3;

assign ap_return_15 = select_ln1495_46_fu_1400_p3;

assign ap_return_16 = select_ln1495_47_fu_1454_p3;

assign ap_return_17 = select_ln1495_48_fu_1508_p3;

assign ap_return_18 = select_ln1495_49_fu_1562_p3;

assign ap_return_19 = select_ln1495_50_fu_1616_p3;

assign ap_return_2 = select_ln1495_33_fu_698_p3;

assign ap_return_20 = select_ln1495_51_fu_1670_p3;

assign ap_return_21 = select_ln1495_52_fu_1724_p3;

assign ap_return_22 = select_ln1495_53_fu_1778_p3;

assign ap_return_23 = select_ln1495_54_fu_1832_p3;

assign ap_return_24 = select_ln1495_55_fu_1886_p3;

assign ap_return_25 = select_ln1495_56_fu_1940_p3;

assign ap_return_26 = select_ln1495_57_fu_1994_p3;

assign ap_return_27 = select_ln1495_58_fu_2048_p3;

assign ap_return_28 = select_ln1495_59_fu_2102_p3;

assign ap_return_29 = select_ln1495_60_fu_2156_p3;

assign ap_return_3 = select_ln1495_34_fu_752_p3;

assign ap_return_30 = select_ln1495_61_fu_2210_p3;

assign ap_return_31 = select_ln1495_62_fu_2264_p3;

assign ap_return_32 = select_ln1495_63_fu_2318_p3;

assign ap_return_33 = select_ln1495_64_fu_2372_p3;

assign ap_return_34 = select_ln1495_65_fu_2426_p3;

assign ap_return_35 = select_ln1495_66_fu_2480_p3;

assign ap_return_36 = select_ln1495_67_fu_2534_p3;

assign ap_return_37 = select_ln1495_68_fu_2588_p3;

assign ap_return_38 = select_ln1495_69_fu_2642_p3;

assign ap_return_39 = select_ln1495_70_fu_2696_p3;

assign ap_return_4 = select_ln1495_35_fu_806_p3;

assign ap_return_40 = select_ln1495_71_fu_2750_p3;

assign ap_return_41 = select_ln1495_72_fu_2804_p3;

assign ap_return_42 = select_ln1495_73_fu_2858_p3;

assign ap_return_43 = select_ln1495_74_fu_2912_p3;

assign ap_return_44 = select_ln1495_75_fu_2966_p3;

assign ap_return_45 = select_ln1495_76_fu_3020_p3;

assign ap_return_46 = select_ln1495_77_fu_3074_p3;

assign ap_return_47 = select_ln1495_78_fu_3128_p3;

assign ap_return_48 = select_ln1495_79_fu_3182_p3;

assign ap_return_49 = select_ln1495_80_fu_3236_p3;

assign ap_return_5 = select_ln1495_36_fu_860_p3;

assign ap_return_50 = select_ln1495_81_fu_3290_p3;

assign ap_return_51 = select_ln1495_82_fu_3344_p3;

assign ap_return_52 = select_ln1495_83_fu_3398_p3;

assign ap_return_53 = select_ln1495_84_fu_3452_p3;

assign ap_return_54 = select_ln1495_85_fu_3506_p3;

assign ap_return_55 = select_ln1495_86_fu_3560_p3;

assign ap_return_56 = select_ln1495_87_fu_3614_p3;

assign ap_return_57 = select_ln1495_88_fu_3668_p3;

assign ap_return_58 = select_ln1495_89_fu_3722_p3;

assign ap_return_59 = select_ln1495_90_fu_3776_p3;

assign ap_return_6 = select_ln1495_37_fu_914_p3;

assign ap_return_60 = select_ln1495_91_fu_3830_p3;

assign ap_return_61 = select_ln1495_92_fu_3884_p3;

assign ap_return_62 = select_ln1495_93_fu_3938_p3;

assign ap_return_63 = select_ln1495_94_fu_3992_p3;

assign ap_return_7 = select_ln1495_38_fu_968_p3;

assign ap_return_8 = select_ln1495_39_fu_1022_p3;

assign ap_return_9 = select_ln1495_40_fu_1076_p3;

assign icmp_ln1494_10_fu_1092_p2 = (((data_10_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_11_fu_1146_p2 = (((data_11_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_12_fu_1200_p2 = (((data_12_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_13_fu_1254_p2 = (((data_13_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_14_fu_1308_p2 = (((data_14_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_15_fu_1362_p2 = (((data_15_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_16_fu_1416_p2 = (((data_16_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_17_fu_1470_p2 = (((data_17_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_18_fu_1524_p2 = (((data_18_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_19_fu_1578_p2 = (((data_19_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_1_fu_606_p2 = (((data_1_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_20_fu_1632_p2 = (((data_20_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_21_fu_1686_p2 = (((data_21_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_22_fu_1740_p2 = (((data_22_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_23_fu_1794_p2 = (((data_23_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_24_fu_1848_p2 = (((data_24_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_25_fu_1902_p2 = (((data_25_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_26_fu_1956_p2 = (((data_26_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_27_fu_2010_p2 = (((data_27_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_28_fu_2064_p2 = (((data_28_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_29_fu_2118_p2 = (((data_29_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_2_fu_660_p2 = (((data_2_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_30_fu_2172_p2 = (((data_30_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_31_fu_2226_p2 = (((data_31_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_32_fu_2280_p2 = (((data_32_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_33_fu_2334_p2 = (((data_33_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_34_fu_2388_p2 = (((data_34_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_35_fu_2442_p2 = (((data_35_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_36_fu_2496_p2 = (((data_36_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_37_fu_2550_p2 = (((data_37_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_38_fu_2604_p2 = (((data_38_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_39_fu_2658_p2 = (((data_39_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_3_fu_714_p2 = (((data_3_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_40_fu_2712_p2 = (((data_40_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_41_fu_2766_p2 = (((data_41_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_42_fu_2820_p2 = (((data_42_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_43_fu_2874_p2 = (((data_43_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_44_fu_2928_p2 = (((data_44_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_45_fu_2982_p2 = (((data_45_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_46_fu_3036_p2 = (((data_46_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_47_fu_3090_p2 = (((data_47_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_48_fu_3144_p2 = (((data_48_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_49_fu_3198_p2 = (((data_49_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_4_fu_768_p2 = (((data_4_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_50_fu_3252_p2 = (((data_50_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_51_fu_3306_p2 = (((data_51_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_52_fu_3360_p2 = (((data_52_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_53_fu_3414_p2 = (((data_53_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_54_fu_3468_p2 = (((data_54_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_55_fu_3522_p2 = (((data_55_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_56_fu_3576_p2 = (((data_56_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_57_fu_3630_p2 = (((data_57_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_58_fu_3684_p2 = (((data_58_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_59_fu_3738_p2 = (((data_59_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_5_fu_822_p2 = (((data_5_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_60_fu_3792_p2 = (((data_60_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_61_fu_3846_p2 = (((data_61_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_62_fu_3900_p2 = (((data_62_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_63_fu_3954_p2 = (((data_63_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_6_fu_876_p2 = (((data_6_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_7_fu_930_p2 = (((data_7_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_8_fu_984_p2 = (((data_8_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_9_fu_1038_p2 = (((data_9_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_fu_552_p2 = (((data_0_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign or_ln1495_32_fu_638_p2 = (tmp_100_fu_598_p3 | icmp_ln1494_1_fu_606_p2);

assign or_ln1495_33_fu_692_p2 = (tmp_103_fu_652_p3 | icmp_ln1494_2_fu_660_p2);

assign or_ln1495_34_fu_746_p2 = (tmp_106_fu_706_p3 | icmp_ln1494_3_fu_714_p2);

assign or_ln1495_35_fu_800_p2 = (tmp_109_fu_760_p3 | icmp_ln1494_4_fu_768_p2);

assign or_ln1495_36_fu_854_p2 = (tmp_112_fu_814_p3 | icmp_ln1494_5_fu_822_p2);

assign or_ln1495_37_fu_908_p2 = (tmp_115_fu_868_p3 | icmp_ln1494_6_fu_876_p2);

assign or_ln1495_38_fu_962_p2 = (tmp_118_fu_922_p3 | icmp_ln1494_7_fu_930_p2);

assign or_ln1495_39_fu_1016_p2 = (tmp_121_fu_976_p3 | icmp_ln1494_8_fu_984_p2);

assign or_ln1495_40_fu_1070_p2 = (tmp_124_fu_1030_p3 | icmp_ln1494_9_fu_1038_p2);

assign or_ln1495_41_fu_1124_p2 = (tmp_127_fu_1084_p3 | icmp_ln1494_10_fu_1092_p2);

assign or_ln1495_42_fu_1178_p2 = (tmp_130_fu_1138_p3 | icmp_ln1494_11_fu_1146_p2);

assign or_ln1495_43_fu_1232_p2 = (tmp_133_fu_1192_p3 | icmp_ln1494_12_fu_1200_p2);

assign or_ln1495_44_fu_1286_p2 = (tmp_136_fu_1246_p3 | icmp_ln1494_13_fu_1254_p2);

assign or_ln1495_45_fu_1340_p2 = (tmp_139_fu_1300_p3 | icmp_ln1494_14_fu_1308_p2);

assign or_ln1495_46_fu_1394_p2 = (tmp_142_fu_1354_p3 | icmp_ln1494_15_fu_1362_p2);

assign or_ln1495_47_fu_1448_p2 = (tmp_145_fu_1408_p3 | icmp_ln1494_16_fu_1416_p2);

assign or_ln1495_48_fu_1502_p2 = (tmp_148_fu_1462_p3 | icmp_ln1494_17_fu_1470_p2);

assign or_ln1495_49_fu_1556_p2 = (tmp_151_fu_1516_p3 | icmp_ln1494_18_fu_1524_p2);

assign or_ln1495_50_fu_1610_p2 = (tmp_154_fu_1570_p3 | icmp_ln1494_19_fu_1578_p2);

assign or_ln1495_51_fu_1664_p2 = (tmp_157_fu_1624_p3 | icmp_ln1494_20_fu_1632_p2);

assign or_ln1495_52_fu_1718_p2 = (tmp_160_fu_1678_p3 | icmp_ln1494_21_fu_1686_p2);

assign or_ln1495_53_fu_1772_p2 = (tmp_163_fu_1732_p3 | icmp_ln1494_22_fu_1740_p2);

assign or_ln1495_54_fu_1826_p2 = (tmp_166_fu_1786_p3 | icmp_ln1494_23_fu_1794_p2);

assign or_ln1495_55_fu_1880_p2 = (tmp_169_fu_1840_p3 | icmp_ln1494_24_fu_1848_p2);

assign or_ln1495_56_fu_1934_p2 = (tmp_172_fu_1894_p3 | icmp_ln1494_25_fu_1902_p2);

assign or_ln1495_57_fu_1988_p2 = (tmp_175_fu_1948_p3 | icmp_ln1494_26_fu_1956_p2);

assign or_ln1495_58_fu_2042_p2 = (tmp_178_fu_2002_p3 | icmp_ln1494_27_fu_2010_p2);

assign or_ln1495_59_fu_2096_p2 = (tmp_181_fu_2056_p3 | icmp_ln1494_28_fu_2064_p2);

assign or_ln1495_60_fu_2150_p2 = (tmp_184_fu_2110_p3 | icmp_ln1494_29_fu_2118_p2);

assign or_ln1495_61_fu_2204_p2 = (tmp_187_fu_2164_p3 | icmp_ln1494_30_fu_2172_p2);

assign or_ln1495_62_fu_2258_p2 = (tmp_190_fu_2218_p3 | icmp_ln1494_31_fu_2226_p2);

assign or_ln1495_63_fu_2312_p2 = (tmp_193_fu_2272_p3 | icmp_ln1494_32_fu_2280_p2);

assign or_ln1495_64_fu_2366_p2 = (tmp_196_fu_2326_p3 | icmp_ln1494_33_fu_2334_p2);

assign or_ln1495_65_fu_2420_p2 = (tmp_199_fu_2380_p3 | icmp_ln1494_34_fu_2388_p2);

assign or_ln1495_66_fu_2474_p2 = (tmp_202_fu_2434_p3 | icmp_ln1494_35_fu_2442_p2);

assign or_ln1495_67_fu_2528_p2 = (tmp_205_fu_2488_p3 | icmp_ln1494_36_fu_2496_p2);

assign or_ln1495_68_fu_2582_p2 = (tmp_208_fu_2542_p3 | icmp_ln1494_37_fu_2550_p2);

assign or_ln1495_69_fu_2636_p2 = (tmp_211_fu_2596_p3 | icmp_ln1494_38_fu_2604_p2);

assign or_ln1495_70_fu_2690_p2 = (tmp_214_fu_2650_p3 | icmp_ln1494_39_fu_2658_p2);

assign or_ln1495_71_fu_2744_p2 = (tmp_217_fu_2704_p3 | icmp_ln1494_40_fu_2712_p2);

assign or_ln1495_72_fu_2798_p2 = (tmp_220_fu_2758_p3 | icmp_ln1494_41_fu_2766_p2);

assign or_ln1495_73_fu_2852_p2 = (tmp_223_fu_2812_p3 | icmp_ln1494_42_fu_2820_p2);

assign or_ln1495_74_fu_2906_p2 = (tmp_226_fu_2866_p3 | icmp_ln1494_43_fu_2874_p2);

assign or_ln1495_75_fu_2960_p2 = (tmp_229_fu_2920_p3 | icmp_ln1494_44_fu_2928_p2);

assign or_ln1495_76_fu_3014_p2 = (tmp_232_fu_2974_p3 | icmp_ln1494_45_fu_2982_p2);

assign or_ln1495_77_fu_3068_p2 = (tmp_235_fu_3028_p3 | icmp_ln1494_46_fu_3036_p2);

assign or_ln1495_78_fu_3122_p2 = (tmp_238_fu_3082_p3 | icmp_ln1494_47_fu_3090_p2);

assign or_ln1495_79_fu_3176_p2 = (tmp_241_fu_3136_p3 | icmp_ln1494_48_fu_3144_p2);

assign or_ln1495_80_fu_3230_p2 = (tmp_244_fu_3190_p3 | icmp_ln1494_49_fu_3198_p2);

assign or_ln1495_81_fu_3284_p2 = (tmp_247_fu_3244_p3 | icmp_ln1494_50_fu_3252_p2);

assign or_ln1495_82_fu_3338_p2 = (tmp_250_fu_3298_p3 | icmp_ln1494_51_fu_3306_p2);

assign or_ln1495_83_fu_3392_p2 = (tmp_253_fu_3352_p3 | icmp_ln1494_52_fu_3360_p2);

assign or_ln1495_84_fu_3446_p2 = (tmp_256_fu_3406_p3 | icmp_ln1494_53_fu_3414_p2);

assign or_ln1495_85_fu_3500_p2 = (tmp_259_fu_3460_p3 | icmp_ln1494_54_fu_3468_p2);

assign or_ln1495_86_fu_3554_p2 = (tmp_262_fu_3514_p3 | icmp_ln1494_55_fu_3522_p2);

assign or_ln1495_87_fu_3608_p2 = (tmp_265_fu_3568_p3 | icmp_ln1494_56_fu_3576_p2);

assign or_ln1495_88_fu_3662_p2 = (tmp_268_fu_3622_p3 | icmp_ln1494_57_fu_3630_p2);

assign or_ln1495_89_fu_3716_p2 = (tmp_271_fu_3676_p3 | icmp_ln1494_58_fu_3684_p2);

assign or_ln1495_90_fu_3770_p2 = (tmp_274_fu_3730_p3 | icmp_ln1494_59_fu_3738_p2);

assign or_ln1495_91_fu_3824_p2 = (tmp_277_fu_3784_p3 | icmp_ln1494_60_fu_3792_p2);

assign or_ln1495_92_fu_3878_p2 = (tmp_280_fu_3838_p3 | icmp_ln1494_61_fu_3846_p2);

assign or_ln1495_93_fu_3932_p2 = (tmp_283_fu_3892_p3 | icmp_ln1494_62_fu_3900_p2);

assign or_ln1495_94_fu_3986_p2 = (tmp_286_fu_3946_p3 | icmp_ln1494_63_fu_3954_p2);

assign or_ln1495_fu_584_p2 = (tmp_97_fu_544_p3 | icmp_ln1494_fu_552_p2);

assign select_ln1495_32_fu_644_p3 = ((or_ln1495_32_fu_638_p2[0:0] == 1'b1) ? zext_ln1495_32_fu_634_p1 : data_1_V_read);

assign select_ln1495_33_fu_698_p3 = ((or_ln1495_33_fu_692_p2[0:0] == 1'b1) ? zext_ln1495_33_fu_688_p1 : data_2_V_read);

assign select_ln1495_34_fu_752_p3 = ((or_ln1495_34_fu_746_p2[0:0] == 1'b1) ? zext_ln1495_34_fu_742_p1 : data_3_V_read);

assign select_ln1495_35_fu_806_p3 = ((or_ln1495_35_fu_800_p2[0:0] == 1'b1) ? zext_ln1495_35_fu_796_p1 : data_4_V_read);

assign select_ln1495_36_fu_860_p3 = ((or_ln1495_36_fu_854_p2[0:0] == 1'b1) ? zext_ln1495_36_fu_850_p1 : data_5_V_read);

assign select_ln1495_37_fu_914_p3 = ((or_ln1495_37_fu_908_p2[0:0] == 1'b1) ? zext_ln1495_37_fu_904_p1 : data_6_V_read);

assign select_ln1495_38_fu_968_p3 = ((or_ln1495_38_fu_962_p2[0:0] == 1'b1) ? zext_ln1495_38_fu_958_p1 : data_7_V_read);

assign select_ln1495_39_fu_1022_p3 = ((or_ln1495_39_fu_1016_p2[0:0] == 1'b1) ? zext_ln1495_39_fu_1012_p1 : data_8_V_read);

assign select_ln1495_40_fu_1076_p3 = ((or_ln1495_40_fu_1070_p2[0:0] == 1'b1) ? zext_ln1495_40_fu_1066_p1 : data_9_V_read);

assign select_ln1495_41_fu_1130_p3 = ((or_ln1495_41_fu_1124_p2[0:0] == 1'b1) ? zext_ln1495_41_fu_1120_p1 : data_10_V_read);

assign select_ln1495_42_fu_1184_p3 = ((or_ln1495_42_fu_1178_p2[0:0] == 1'b1) ? zext_ln1495_42_fu_1174_p1 : data_11_V_read);

assign select_ln1495_43_fu_1238_p3 = ((or_ln1495_43_fu_1232_p2[0:0] == 1'b1) ? zext_ln1495_43_fu_1228_p1 : data_12_V_read);

assign select_ln1495_44_fu_1292_p3 = ((or_ln1495_44_fu_1286_p2[0:0] == 1'b1) ? zext_ln1495_44_fu_1282_p1 : data_13_V_read);

assign select_ln1495_45_fu_1346_p3 = ((or_ln1495_45_fu_1340_p2[0:0] == 1'b1) ? zext_ln1495_45_fu_1336_p1 : data_14_V_read);

assign select_ln1495_46_fu_1400_p3 = ((or_ln1495_46_fu_1394_p2[0:0] == 1'b1) ? zext_ln1495_46_fu_1390_p1 : data_15_V_read);

assign select_ln1495_47_fu_1454_p3 = ((or_ln1495_47_fu_1448_p2[0:0] == 1'b1) ? zext_ln1495_47_fu_1444_p1 : data_16_V_read);

assign select_ln1495_48_fu_1508_p3 = ((or_ln1495_48_fu_1502_p2[0:0] == 1'b1) ? zext_ln1495_48_fu_1498_p1 : data_17_V_read);

assign select_ln1495_49_fu_1562_p3 = ((or_ln1495_49_fu_1556_p2[0:0] == 1'b1) ? zext_ln1495_49_fu_1552_p1 : data_18_V_read);

assign select_ln1495_50_fu_1616_p3 = ((or_ln1495_50_fu_1610_p2[0:0] == 1'b1) ? zext_ln1495_50_fu_1606_p1 : data_19_V_read);

assign select_ln1495_51_fu_1670_p3 = ((or_ln1495_51_fu_1664_p2[0:0] == 1'b1) ? zext_ln1495_51_fu_1660_p1 : data_20_V_read);

assign select_ln1495_52_fu_1724_p3 = ((or_ln1495_52_fu_1718_p2[0:0] == 1'b1) ? zext_ln1495_52_fu_1714_p1 : data_21_V_read);

assign select_ln1495_53_fu_1778_p3 = ((or_ln1495_53_fu_1772_p2[0:0] == 1'b1) ? zext_ln1495_53_fu_1768_p1 : data_22_V_read);

assign select_ln1495_54_fu_1832_p3 = ((or_ln1495_54_fu_1826_p2[0:0] == 1'b1) ? zext_ln1495_54_fu_1822_p1 : data_23_V_read);

assign select_ln1495_55_fu_1886_p3 = ((or_ln1495_55_fu_1880_p2[0:0] == 1'b1) ? zext_ln1495_55_fu_1876_p1 : data_24_V_read);

assign select_ln1495_56_fu_1940_p3 = ((or_ln1495_56_fu_1934_p2[0:0] == 1'b1) ? zext_ln1495_56_fu_1930_p1 : data_25_V_read);

assign select_ln1495_57_fu_1994_p3 = ((or_ln1495_57_fu_1988_p2[0:0] == 1'b1) ? zext_ln1495_57_fu_1984_p1 : data_26_V_read);

assign select_ln1495_58_fu_2048_p3 = ((or_ln1495_58_fu_2042_p2[0:0] == 1'b1) ? zext_ln1495_58_fu_2038_p1 : data_27_V_read);

assign select_ln1495_59_fu_2102_p3 = ((or_ln1495_59_fu_2096_p2[0:0] == 1'b1) ? zext_ln1495_59_fu_2092_p1 : data_28_V_read);

assign select_ln1495_60_fu_2156_p3 = ((or_ln1495_60_fu_2150_p2[0:0] == 1'b1) ? zext_ln1495_60_fu_2146_p1 : data_29_V_read);

assign select_ln1495_61_fu_2210_p3 = ((or_ln1495_61_fu_2204_p2[0:0] == 1'b1) ? zext_ln1495_61_fu_2200_p1 : data_30_V_read);

assign select_ln1495_62_fu_2264_p3 = ((or_ln1495_62_fu_2258_p2[0:0] == 1'b1) ? zext_ln1495_62_fu_2254_p1 : data_31_V_read);

assign select_ln1495_63_fu_2318_p3 = ((or_ln1495_63_fu_2312_p2[0:0] == 1'b1) ? zext_ln1495_63_fu_2308_p1 : data_32_V_read);

assign select_ln1495_64_fu_2372_p3 = ((or_ln1495_64_fu_2366_p2[0:0] == 1'b1) ? zext_ln1495_64_fu_2362_p1 : data_33_V_read);

assign select_ln1495_65_fu_2426_p3 = ((or_ln1495_65_fu_2420_p2[0:0] == 1'b1) ? zext_ln1495_65_fu_2416_p1 : data_34_V_read);

assign select_ln1495_66_fu_2480_p3 = ((or_ln1495_66_fu_2474_p2[0:0] == 1'b1) ? zext_ln1495_66_fu_2470_p1 : data_35_V_read);

assign select_ln1495_67_fu_2534_p3 = ((or_ln1495_67_fu_2528_p2[0:0] == 1'b1) ? zext_ln1495_67_fu_2524_p1 : data_36_V_read);

assign select_ln1495_68_fu_2588_p3 = ((or_ln1495_68_fu_2582_p2[0:0] == 1'b1) ? zext_ln1495_68_fu_2578_p1 : data_37_V_read);

assign select_ln1495_69_fu_2642_p3 = ((or_ln1495_69_fu_2636_p2[0:0] == 1'b1) ? zext_ln1495_69_fu_2632_p1 : data_38_V_read);

assign select_ln1495_70_fu_2696_p3 = ((or_ln1495_70_fu_2690_p2[0:0] == 1'b1) ? zext_ln1495_70_fu_2686_p1 : data_39_V_read);

assign select_ln1495_71_fu_2750_p3 = ((or_ln1495_71_fu_2744_p2[0:0] == 1'b1) ? zext_ln1495_71_fu_2740_p1 : data_40_V_read);

assign select_ln1495_72_fu_2804_p3 = ((or_ln1495_72_fu_2798_p2[0:0] == 1'b1) ? zext_ln1495_72_fu_2794_p1 : data_41_V_read);

assign select_ln1495_73_fu_2858_p3 = ((or_ln1495_73_fu_2852_p2[0:0] == 1'b1) ? zext_ln1495_73_fu_2848_p1 : data_42_V_read);

assign select_ln1495_74_fu_2912_p3 = ((or_ln1495_74_fu_2906_p2[0:0] == 1'b1) ? zext_ln1495_74_fu_2902_p1 : data_43_V_read);

assign select_ln1495_75_fu_2966_p3 = ((or_ln1495_75_fu_2960_p2[0:0] == 1'b1) ? zext_ln1495_75_fu_2956_p1 : data_44_V_read);

assign select_ln1495_76_fu_3020_p3 = ((or_ln1495_76_fu_3014_p2[0:0] == 1'b1) ? zext_ln1495_76_fu_3010_p1 : data_45_V_read);

assign select_ln1495_77_fu_3074_p3 = ((or_ln1495_77_fu_3068_p2[0:0] == 1'b1) ? zext_ln1495_77_fu_3064_p1 : data_46_V_read);

assign select_ln1495_78_fu_3128_p3 = ((or_ln1495_78_fu_3122_p2[0:0] == 1'b1) ? zext_ln1495_78_fu_3118_p1 : data_47_V_read);

assign select_ln1495_79_fu_3182_p3 = ((or_ln1495_79_fu_3176_p2[0:0] == 1'b1) ? zext_ln1495_79_fu_3172_p1 : data_48_V_read);

assign select_ln1495_80_fu_3236_p3 = ((or_ln1495_80_fu_3230_p2[0:0] == 1'b1) ? zext_ln1495_80_fu_3226_p1 : data_49_V_read);

assign select_ln1495_81_fu_3290_p3 = ((or_ln1495_81_fu_3284_p2[0:0] == 1'b1) ? zext_ln1495_81_fu_3280_p1 : data_50_V_read);

assign select_ln1495_82_fu_3344_p3 = ((or_ln1495_82_fu_3338_p2[0:0] == 1'b1) ? zext_ln1495_82_fu_3334_p1 : data_51_V_read);

assign select_ln1495_83_fu_3398_p3 = ((or_ln1495_83_fu_3392_p2[0:0] == 1'b1) ? zext_ln1495_83_fu_3388_p1 : data_52_V_read);

assign select_ln1495_84_fu_3452_p3 = ((or_ln1495_84_fu_3446_p2[0:0] == 1'b1) ? zext_ln1495_84_fu_3442_p1 : data_53_V_read);

assign select_ln1495_85_fu_3506_p3 = ((or_ln1495_85_fu_3500_p2[0:0] == 1'b1) ? zext_ln1495_85_fu_3496_p1 : data_54_V_read);

assign select_ln1495_86_fu_3560_p3 = ((or_ln1495_86_fu_3554_p2[0:0] == 1'b1) ? zext_ln1495_86_fu_3550_p1 : data_55_V_read);

assign select_ln1495_87_fu_3614_p3 = ((or_ln1495_87_fu_3608_p2[0:0] == 1'b1) ? zext_ln1495_87_fu_3604_p1 : data_56_V_read);

assign select_ln1495_88_fu_3668_p3 = ((or_ln1495_88_fu_3662_p2[0:0] == 1'b1) ? zext_ln1495_88_fu_3658_p1 : data_57_V_read);

assign select_ln1495_89_fu_3722_p3 = ((or_ln1495_89_fu_3716_p2[0:0] == 1'b1) ? zext_ln1495_89_fu_3712_p1 : data_58_V_read);

assign select_ln1495_90_fu_3776_p3 = ((or_ln1495_90_fu_3770_p2[0:0] == 1'b1) ? zext_ln1495_90_fu_3766_p1 : data_59_V_read);

assign select_ln1495_91_fu_3830_p3 = ((or_ln1495_91_fu_3824_p2[0:0] == 1'b1) ? zext_ln1495_91_fu_3820_p1 : data_60_V_read);

assign select_ln1495_92_fu_3884_p3 = ((or_ln1495_92_fu_3878_p2[0:0] == 1'b1) ? zext_ln1495_92_fu_3874_p1 : data_61_V_read);

assign select_ln1495_93_fu_3938_p3 = ((or_ln1495_93_fu_3932_p2[0:0] == 1'b1) ? zext_ln1495_93_fu_3928_p1 : data_62_V_read);

assign select_ln1495_94_fu_3992_p3 = ((or_ln1495_94_fu_3986_p2[0:0] == 1'b1) ? zext_ln1495_94_fu_3982_p1 : data_63_V_read);

assign select_ln1495_fu_590_p3 = ((or_ln1495_fu_584_p2[0:0] == 1'b1) ? zext_ln1495_fu_580_p1 : data_0_V_read);

assign tmp_100_fu_598_p3 = data_1_V_read[32'd15];

assign tmp_101_fu_612_p3 = data_1_V_read[32'd15];

assign tmp_102_fu_626_p3 = {{xor_ln1495_32_fu_620_p2}, {10'd0}};

assign tmp_103_fu_652_p3 = data_2_V_read[32'd15];

assign tmp_104_fu_666_p3 = data_2_V_read[32'd15];

assign tmp_105_fu_680_p3 = {{xor_ln1495_33_fu_674_p2}, {10'd0}};

assign tmp_106_fu_706_p3 = data_3_V_read[32'd15];

assign tmp_107_fu_720_p3 = data_3_V_read[32'd15];

assign tmp_108_fu_734_p3 = {{xor_ln1495_34_fu_728_p2}, {10'd0}};

assign tmp_109_fu_760_p3 = data_4_V_read[32'd15];

assign tmp_110_fu_774_p3 = data_4_V_read[32'd15];

assign tmp_111_fu_788_p3 = {{xor_ln1495_35_fu_782_p2}, {10'd0}};

assign tmp_112_fu_814_p3 = data_5_V_read[32'd15];

assign tmp_113_fu_828_p3 = data_5_V_read[32'd15];

assign tmp_114_fu_842_p3 = {{xor_ln1495_36_fu_836_p2}, {10'd0}};

assign tmp_115_fu_868_p3 = data_6_V_read[32'd15];

assign tmp_116_fu_882_p3 = data_6_V_read[32'd15];

assign tmp_117_fu_896_p3 = {{xor_ln1495_37_fu_890_p2}, {10'd0}};

assign tmp_118_fu_922_p3 = data_7_V_read[32'd15];

assign tmp_119_fu_936_p3 = data_7_V_read[32'd15];

assign tmp_120_fu_950_p3 = {{xor_ln1495_38_fu_944_p2}, {10'd0}};

assign tmp_121_fu_976_p3 = data_8_V_read[32'd15];

assign tmp_122_fu_990_p3 = data_8_V_read[32'd15];

assign tmp_123_fu_1004_p3 = {{xor_ln1495_39_fu_998_p2}, {10'd0}};

assign tmp_124_fu_1030_p3 = data_9_V_read[32'd15];

assign tmp_125_fu_1044_p3 = data_9_V_read[32'd15];

assign tmp_126_fu_1058_p3 = {{xor_ln1495_40_fu_1052_p2}, {10'd0}};

assign tmp_127_fu_1084_p3 = data_10_V_read[32'd15];

assign tmp_128_fu_1098_p3 = data_10_V_read[32'd15];

assign tmp_129_fu_1112_p3 = {{xor_ln1495_41_fu_1106_p2}, {10'd0}};

assign tmp_130_fu_1138_p3 = data_11_V_read[32'd15];

assign tmp_131_fu_1152_p3 = data_11_V_read[32'd15];

assign tmp_132_fu_1166_p3 = {{xor_ln1495_42_fu_1160_p2}, {10'd0}};

assign tmp_133_fu_1192_p3 = data_12_V_read[32'd15];

assign tmp_134_fu_1206_p3 = data_12_V_read[32'd15];

assign tmp_135_fu_1220_p3 = {{xor_ln1495_43_fu_1214_p2}, {10'd0}};

assign tmp_136_fu_1246_p3 = data_13_V_read[32'd15];

assign tmp_137_fu_1260_p3 = data_13_V_read[32'd15];

assign tmp_138_fu_1274_p3 = {{xor_ln1495_44_fu_1268_p2}, {10'd0}};

assign tmp_139_fu_1300_p3 = data_14_V_read[32'd15];

assign tmp_140_fu_1314_p3 = data_14_V_read[32'd15];

assign tmp_141_fu_1328_p3 = {{xor_ln1495_45_fu_1322_p2}, {10'd0}};

assign tmp_142_fu_1354_p3 = data_15_V_read[32'd15];

assign tmp_143_fu_1368_p3 = data_15_V_read[32'd15];

assign tmp_144_fu_1382_p3 = {{xor_ln1495_46_fu_1376_p2}, {10'd0}};

assign tmp_145_fu_1408_p3 = data_16_V_read[32'd15];

assign tmp_146_fu_1422_p3 = data_16_V_read[32'd15];

assign tmp_147_fu_1436_p3 = {{xor_ln1495_47_fu_1430_p2}, {10'd0}};

assign tmp_148_fu_1462_p3 = data_17_V_read[32'd15];

assign tmp_149_fu_1476_p3 = data_17_V_read[32'd15];

assign tmp_150_fu_1490_p3 = {{xor_ln1495_48_fu_1484_p2}, {10'd0}};

assign tmp_151_fu_1516_p3 = data_18_V_read[32'd15];

assign tmp_152_fu_1530_p3 = data_18_V_read[32'd15];

assign tmp_153_fu_1544_p3 = {{xor_ln1495_49_fu_1538_p2}, {10'd0}};

assign tmp_154_fu_1570_p3 = data_19_V_read[32'd15];

assign tmp_155_fu_1584_p3 = data_19_V_read[32'd15];

assign tmp_156_fu_1598_p3 = {{xor_ln1495_50_fu_1592_p2}, {10'd0}};

assign tmp_157_fu_1624_p3 = data_20_V_read[32'd15];

assign tmp_158_fu_1638_p3 = data_20_V_read[32'd15];

assign tmp_159_fu_1652_p3 = {{xor_ln1495_51_fu_1646_p2}, {10'd0}};

assign tmp_160_fu_1678_p3 = data_21_V_read[32'd15];

assign tmp_161_fu_1692_p3 = data_21_V_read[32'd15];

assign tmp_162_fu_1706_p3 = {{xor_ln1495_52_fu_1700_p2}, {10'd0}};

assign tmp_163_fu_1732_p3 = data_22_V_read[32'd15];

assign tmp_164_fu_1746_p3 = data_22_V_read[32'd15];

assign tmp_165_fu_1760_p3 = {{xor_ln1495_53_fu_1754_p2}, {10'd0}};

assign tmp_166_fu_1786_p3 = data_23_V_read[32'd15];

assign tmp_167_fu_1800_p3 = data_23_V_read[32'd15];

assign tmp_168_fu_1814_p3 = {{xor_ln1495_54_fu_1808_p2}, {10'd0}};

assign tmp_169_fu_1840_p3 = data_24_V_read[32'd15];

assign tmp_170_fu_1854_p3 = data_24_V_read[32'd15];

assign tmp_171_fu_1868_p3 = {{xor_ln1495_55_fu_1862_p2}, {10'd0}};

assign tmp_172_fu_1894_p3 = data_25_V_read[32'd15];

assign tmp_173_fu_1908_p3 = data_25_V_read[32'd15];

assign tmp_174_fu_1922_p3 = {{xor_ln1495_56_fu_1916_p2}, {10'd0}};

assign tmp_175_fu_1948_p3 = data_26_V_read[32'd15];

assign tmp_176_fu_1962_p3 = data_26_V_read[32'd15];

assign tmp_177_fu_1976_p3 = {{xor_ln1495_57_fu_1970_p2}, {10'd0}};

assign tmp_178_fu_2002_p3 = data_27_V_read[32'd15];

assign tmp_179_fu_2016_p3 = data_27_V_read[32'd15];

assign tmp_180_fu_2030_p3 = {{xor_ln1495_58_fu_2024_p2}, {10'd0}};

assign tmp_181_fu_2056_p3 = data_28_V_read[32'd15];

assign tmp_182_fu_2070_p3 = data_28_V_read[32'd15];

assign tmp_183_fu_2084_p3 = {{xor_ln1495_59_fu_2078_p2}, {10'd0}};

assign tmp_184_fu_2110_p3 = data_29_V_read[32'd15];

assign tmp_185_fu_2124_p3 = data_29_V_read[32'd15];

assign tmp_186_fu_2138_p3 = {{xor_ln1495_60_fu_2132_p2}, {10'd0}};

assign tmp_187_fu_2164_p3 = data_30_V_read[32'd15];

assign tmp_188_fu_2178_p3 = data_30_V_read[32'd15];

assign tmp_189_fu_2192_p3 = {{xor_ln1495_61_fu_2186_p2}, {10'd0}};

assign tmp_190_fu_2218_p3 = data_31_V_read[32'd15];

assign tmp_191_fu_2232_p3 = data_31_V_read[32'd15];

assign tmp_192_fu_2246_p3 = {{xor_ln1495_62_fu_2240_p2}, {10'd0}};

assign tmp_193_fu_2272_p3 = data_32_V_read[32'd15];

assign tmp_194_fu_2286_p3 = data_32_V_read[32'd15];

assign tmp_195_fu_2300_p3 = {{xor_ln1495_63_fu_2294_p2}, {10'd0}};

assign tmp_196_fu_2326_p3 = data_33_V_read[32'd15];

assign tmp_197_fu_2340_p3 = data_33_V_read[32'd15];

assign tmp_198_fu_2354_p3 = {{xor_ln1495_64_fu_2348_p2}, {10'd0}};

assign tmp_199_fu_2380_p3 = data_34_V_read[32'd15];

assign tmp_200_fu_2394_p3 = data_34_V_read[32'd15];

assign tmp_201_fu_2408_p3 = {{xor_ln1495_65_fu_2402_p2}, {10'd0}};

assign tmp_202_fu_2434_p3 = data_35_V_read[32'd15];

assign tmp_203_fu_2448_p3 = data_35_V_read[32'd15];

assign tmp_204_fu_2462_p3 = {{xor_ln1495_66_fu_2456_p2}, {10'd0}};

assign tmp_205_fu_2488_p3 = data_36_V_read[32'd15];

assign tmp_206_fu_2502_p3 = data_36_V_read[32'd15];

assign tmp_207_fu_2516_p3 = {{xor_ln1495_67_fu_2510_p2}, {10'd0}};

assign tmp_208_fu_2542_p3 = data_37_V_read[32'd15];

assign tmp_209_fu_2556_p3 = data_37_V_read[32'd15];

assign tmp_210_fu_2570_p3 = {{xor_ln1495_68_fu_2564_p2}, {10'd0}};

assign tmp_211_fu_2596_p3 = data_38_V_read[32'd15];

assign tmp_212_fu_2610_p3 = data_38_V_read[32'd15];

assign tmp_213_fu_2624_p3 = {{xor_ln1495_69_fu_2618_p2}, {10'd0}};

assign tmp_214_fu_2650_p3 = data_39_V_read[32'd15];

assign tmp_215_fu_2664_p3 = data_39_V_read[32'd15];

assign tmp_216_fu_2678_p3 = {{xor_ln1495_70_fu_2672_p2}, {10'd0}};

assign tmp_217_fu_2704_p3 = data_40_V_read[32'd15];

assign tmp_218_fu_2718_p3 = data_40_V_read[32'd15];

assign tmp_219_fu_2732_p3 = {{xor_ln1495_71_fu_2726_p2}, {10'd0}};

assign tmp_220_fu_2758_p3 = data_41_V_read[32'd15];

assign tmp_221_fu_2772_p3 = data_41_V_read[32'd15];

assign tmp_222_fu_2786_p3 = {{xor_ln1495_72_fu_2780_p2}, {10'd0}};

assign tmp_223_fu_2812_p3 = data_42_V_read[32'd15];

assign tmp_224_fu_2826_p3 = data_42_V_read[32'd15];

assign tmp_225_fu_2840_p3 = {{xor_ln1495_73_fu_2834_p2}, {10'd0}};

assign tmp_226_fu_2866_p3 = data_43_V_read[32'd15];

assign tmp_227_fu_2880_p3 = data_43_V_read[32'd15];

assign tmp_228_fu_2894_p3 = {{xor_ln1495_74_fu_2888_p2}, {10'd0}};

assign tmp_229_fu_2920_p3 = data_44_V_read[32'd15];

assign tmp_230_fu_2934_p3 = data_44_V_read[32'd15];

assign tmp_231_fu_2948_p3 = {{xor_ln1495_75_fu_2942_p2}, {10'd0}};

assign tmp_232_fu_2974_p3 = data_45_V_read[32'd15];

assign tmp_233_fu_2988_p3 = data_45_V_read[32'd15];

assign tmp_234_fu_3002_p3 = {{xor_ln1495_76_fu_2996_p2}, {10'd0}};

assign tmp_235_fu_3028_p3 = data_46_V_read[32'd15];

assign tmp_236_fu_3042_p3 = data_46_V_read[32'd15];

assign tmp_237_fu_3056_p3 = {{xor_ln1495_77_fu_3050_p2}, {10'd0}};

assign tmp_238_fu_3082_p3 = data_47_V_read[32'd15];

assign tmp_239_fu_3096_p3 = data_47_V_read[32'd15];

assign tmp_240_fu_3110_p3 = {{xor_ln1495_78_fu_3104_p2}, {10'd0}};

assign tmp_241_fu_3136_p3 = data_48_V_read[32'd15];

assign tmp_242_fu_3150_p3 = data_48_V_read[32'd15];

assign tmp_243_fu_3164_p3 = {{xor_ln1495_79_fu_3158_p2}, {10'd0}};

assign tmp_244_fu_3190_p3 = data_49_V_read[32'd15];

assign tmp_245_fu_3204_p3 = data_49_V_read[32'd15];

assign tmp_246_fu_3218_p3 = {{xor_ln1495_80_fu_3212_p2}, {10'd0}};

assign tmp_247_fu_3244_p3 = data_50_V_read[32'd15];

assign tmp_248_fu_3258_p3 = data_50_V_read[32'd15];

assign tmp_249_fu_3272_p3 = {{xor_ln1495_81_fu_3266_p2}, {10'd0}};

assign tmp_250_fu_3298_p3 = data_51_V_read[32'd15];

assign tmp_251_fu_3312_p3 = data_51_V_read[32'd15];

assign tmp_252_fu_3326_p3 = {{xor_ln1495_82_fu_3320_p2}, {10'd0}};

assign tmp_253_fu_3352_p3 = data_52_V_read[32'd15];

assign tmp_254_fu_3366_p3 = data_52_V_read[32'd15];

assign tmp_255_fu_3380_p3 = {{xor_ln1495_83_fu_3374_p2}, {10'd0}};

assign tmp_256_fu_3406_p3 = data_53_V_read[32'd15];

assign tmp_257_fu_3420_p3 = data_53_V_read[32'd15];

assign tmp_258_fu_3434_p3 = {{xor_ln1495_84_fu_3428_p2}, {10'd0}};

assign tmp_259_fu_3460_p3 = data_54_V_read[32'd15];

assign tmp_260_fu_3474_p3 = data_54_V_read[32'd15];

assign tmp_261_fu_3488_p3 = {{xor_ln1495_85_fu_3482_p2}, {10'd0}};

assign tmp_262_fu_3514_p3 = data_55_V_read[32'd15];

assign tmp_263_fu_3528_p3 = data_55_V_read[32'd15];

assign tmp_264_fu_3542_p3 = {{xor_ln1495_86_fu_3536_p2}, {10'd0}};

assign tmp_265_fu_3568_p3 = data_56_V_read[32'd15];

assign tmp_266_fu_3582_p3 = data_56_V_read[32'd15];

assign tmp_267_fu_3596_p3 = {{xor_ln1495_87_fu_3590_p2}, {10'd0}};

assign tmp_268_fu_3622_p3 = data_57_V_read[32'd15];

assign tmp_269_fu_3636_p3 = data_57_V_read[32'd15];

assign tmp_270_fu_3650_p3 = {{xor_ln1495_88_fu_3644_p2}, {10'd0}};

assign tmp_271_fu_3676_p3 = data_58_V_read[32'd15];

assign tmp_272_fu_3690_p3 = data_58_V_read[32'd15];

assign tmp_273_fu_3704_p3 = {{xor_ln1495_89_fu_3698_p2}, {10'd0}};

assign tmp_274_fu_3730_p3 = data_59_V_read[32'd15];

assign tmp_275_fu_3744_p3 = data_59_V_read[32'd15];

assign tmp_276_fu_3758_p3 = {{xor_ln1495_90_fu_3752_p2}, {10'd0}};

assign tmp_277_fu_3784_p3 = data_60_V_read[32'd15];

assign tmp_278_fu_3798_p3 = data_60_V_read[32'd15];

assign tmp_279_fu_3812_p3 = {{xor_ln1495_91_fu_3806_p2}, {10'd0}};

assign tmp_280_fu_3838_p3 = data_61_V_read[32'd15];

assign tmp_281_fu_3852_p3 = data_61_V_read[32'd15];

assign tmp_282_fu_3866_p3 = {{xor_ln1495_92_fu_3860_p2}, {10'd0}};

assign tmp_283_fu_3892_p3 = data_62_V_read[32'd15];

assign tmp_284_fu_3906_p3 = data_62_V_read[32'd15];

assign tmp_285_fu_3920_p3 = {{xor_ln1495_93_fu_3914_p2}, {10'd0}};

assign tmp_286_fu_3946_p3 = data_63_V_read[32'd15];

assign tmp_287_fu_3960_p3 = data_63_V_read[32'd15];

assign tmp_288_fu_3974_p3 = {{xor_ln1495_94_fu_3968_p2}, {10'd0}};

assign tmp_97_fu_544_p3 = data_0_V_read[32'd15];

assign tmp_98_fu_558_p3 = data_0_V_read[32'd15];

assign tmp_99_fu_572_p3 = {{xor_ln1495_fu_566_p2}, {10'd0}};

assign xor_ln1495_32_fu_620_p2 = (tmp_101_fu_612_p3 ^ 1'd1);

assign xor_ln1495_33_fu_674_p2 = (tmp_104_fu_666_p3 ^ 1'd1);

assign xor_ln1495_34_fu_728_p2 = (tmp_107_fu_720_p3 ^ 1'd1);

assign xor_ln1495_35_fu_782_p2 = (tmp_110_fu_774_p3 ^ 1'd1);

assign xor_ln1495_36_fu_836_p2 = (tmp_113_fu_828_p3 ^ 1'd1);

assign xor_ln1495_37_fu_890_p2 = (tmp_116_fu_882_p3 ^ 1'd1);

assign xor_ln1495_38_fu_944_p2 = (tmp_119_fu_936_p3 ^ 1'd1);

assign xor_ln1495_39_fu_998_p2 = (tmp_122_fu_990_p3 ^ 1'd1);

assign xor_ln1495_40_fu_1052_p2 = (tmp_125_fu_1044_p3 ^ 1'd1);

assign xor_ln1495_41_fu_1106_p2 = (tmp_128_fu_1098_p3 ^ 1'd1);

assign xor_ln1495_42_fu_1160_p2 = (tmp_131_fu_1152_p3 ^ 1'd1);

assign xor_ln1495_43_fu_1214_p2 = (tmp_134_fu_1206_p3 ^ 1'd1);

assign xor_ln1495_44_fu_1268_p2 = (tmp_137_fu_1260_p3 ^ 1'd1);

assign xor_ln1495_45_fu_1322_p2 = (tmp_140_fu_1314_p3 ^ 1'd1);

assign xor_ln1495_46_fu_1376_p2 = (tmp_143_fu_1368_p3 ^ 1'd1);

assign xor_ln1495_47_fu_1430_p2 = (tmp_146_fu_1422_p3 ^ 1'd1);

assign xor_ln1495_48_fu_1484_p2 = (tmp_149_fu_1476_p3 ^ 1'd1);

assign xor_ln1495_49_fu_1538_p2 = (tmp_152_fu_1530_p3 ^ 1'd1);

assign xor_ln1495_50_fu_1592_p2 = (tmp_155_fu_1584_p3 ^ 1'd1);

assign xor_ln1495_51_fu_1646_p2 = (tmp_158_fu_1638_p3 ^ 1'd1);

assign xor_ln1495_52_fu_1700_p2 = (tmp_161_fu_1692_p3 ^ 1'd1);

assign xor_ln1495_53_fu_1754_p2 = (tmp_164_fu_1746_p3 ^ 1'd1);

assign xor_ln1495_54_fu_1808_p2 = (tmp_167_fu_1800_p3 ^ 1'd1);

assign xor_ln1495_55_fu_1862_p2 = (tmp_170_fu_1854_p3 ^ 1'd1);

assign xor_ln1495_56_fu_1916_p2 = (tmp_173_fu_1908_p3 ^ 1'd1);

assign xor_ln1495_57_fu_1970_p2 = (tmp_176_fu_1962_p3 ^ 1'd1);

assign xor_ln1495_58_fu_2024_p2 = (tmp_179_fu_2016_p3 ^ 1'd1);

assign xor_ln1495_59_fu_2078_p2 = (tmp_182_fu_2070_p3 ^ 1'd1);

assign xor_ln1495_60_fu_2132_p2 = (tmp_185_fu_2124_p3 ^ 1'd1);

assign xor_ln1495_61_fu_2186_p2 = (tmp_188_fu_2178_p3 ^ 1'd1);

assign xor_ln1495_62_fu_2240_p2 = (tmp_191_fu_2232_p3 ^ 1'd1);

assign xor_ln1495_63_fu_2294_p2 = (tmp_194_fu_2286_p3 ^ 1'd1);

assign xor_ln1495_64_fu_2348_p2 = (tmp_197_fu_2340_p3 ^ 1'd1);

assign xor_ln1495_65_fu_2402_p2 = (tmp_200_fu_2394_p3 ^ 1'd1);

assign xor_ln1495_66_fu_2456_p2 = (tmp_203_fu_2448_p3 ^ 1'd1);

assign xor_ln1495_67_fu_2510_p2 = (tmp_206_fu_2502_p3 ^ 1'd1);

assign xor_ln1495_68_fu_2564_p2 = (tmp_209_fu_2556_p3 ^ 1'd1);

assign xor_ln1495_69_fu_2618_p2 = (tmp_212_fu_2610_p3 ^ 1'd1);

assign xor_ln1495_70_fu_2672_p2 = (tmp_215_fu_2664_p3 ^ 1'd1);

assign xor_ln1495_71_fu_2726_p2 = (tmp_218_fu_2718_p3 ^ 1'd1);

assign xor_ln1495_72_fu_2780_p2 = (tmp_221_fu_2772_p3 ^ 1'd1);

assign xor_ln1495_73_fu_2834_p2 = (tmp_224_fu_2826_p3 ^ 1'd1);

assign xor_ln1495_74_fu_2888_p2 = (tmp_227_fu_2880_p3 ^ 1'd1);

assign xor_ln1495_75_fu_2942_p2 = (tmp_230_fu_2934_p3 ^ 1'd1);

assign xor_ln1495_76_fu_2996_p2 = (tmp_233_fu_2988_p3 ^ 1'd1);

assign xor_ln1495_77_fu_3050_p2 = (tmp_236_fu_3042_p3 ^ 1'd1);

assign xor_ln1495_78_fu_3104_p2 = (tmp_239_fu_3096_p3 ^ 1'd1);

assign xor_ln1495_79_fu_3158_p2 = (tmp_242_fu_3150_p3 ^ 1'd1);

assign xor_ln1495_80_fu_3212_p2 = (tmp_245_fu_3204_p3 ^ 1'd1);

assign xor_ln1495_81_fu_3266_p2 = (tmp_248_fu_3258_p3 ^ 1'd1);

assign xor_ln1495_82_fu_3320_p2 = (tmp_251_fu_3312_p3 ^ 1'd1);

assign xor_ln1495_83_fu_3374_p2 = (tmp_254_fu_3366_p3 ^ 1'd1);

assign xor_ln1495_84_fu_3428_p2 = (tmp_257_fu_3420_p3 ^ 1'd1);

assign xor_ln1495_85_fu_3482_p2 = (tmp_260_fu_3474_p3 ^ 1'd1);

assign xor_ln1495_86_fu_3536_p2 = (tmp_263_fu_3528_p3 ^ 1'd1);

assign xor_ln1495_87_fu_3590_p2 = (tmp_266_fu_3582_p3 ^ 1'd1);

assign xor_ln1495_88_fu_3644_p2 = (tmp_269_fu_3636_p3 ^ 1'd1);

assign xor_ln1495_89_fu_3698_p2 = (tmp_272_fu_3690_p3 ^ 1'd1);

assign xor_ln1495_90_fu_3752_p2 = (tmp_275_fu_3744_p3 ^ 1'd1);

assign xor_ln1495_91_fu_3806_p2 = (tmp_278_fu_3798_p3 ^ 1'd1);

assign xor_ln1495_92_fu_3860_p2 = (tmp_281_fu_3852_p3 ^ 1'd1);

assign xor_ln1495_93_fu_3914_p2 = (tmp_284_fu_3906_p3 ^ 1'd1);

assign xor_ln1495_94_fu_3968_p2 = (tmp_287_fu_3960_p3 ^ 1'd1);

assign xor_ln1495_fu_566_p2 = (tmp_98_fu_558_p3 ^ 1'd1);

assign zext_ln1495_32_fu_634_p1 = tmp_102_fu_626_p3;

assign zext_ln1495_33_fu_688_p1 = tmp_105_fu_680_p3;

assign zext_ln1495_34_fu_742_p1 = tmp_108_fu_734_p3;

assign zext_ln1495_35_fu_796_p1 = tmp_111_fu_788_p3;

assign zext_ln1495_36_fu_850_p1 = tmp_114_fu_842_p3;

assign zext_ln1495_37_fu_904_p1 = tmp_117_fu_896_p3;

assign zext_ln1495_38_fu_958_p1 = tmp_120_fu_950_p3;

assign zext_ln1495_39_fu_1012_p1 = tmp_123_fu_1004_p3;

assign zext_ln1495_40_fu_1066_p1 = tmp_126_fu_1058_p3;

assign zext_ln1495_41_fu_1120_p1 = tmp_129_fu_1112_p3;

assign zext_ln1495_42_fu_1174_p1 = tmp_132_fu_1166_p3;

assign zext_ln1495_43_fu_1228_p1 = tmp_135_fu_1220_p3;

assign zext_ln1495_44_fu_1282_p1 = tmp_138_fu_1274_p3;

assign zext_ln1495_45_fu_1336_p1 = tmp_141_fu_1328_p3;

assign zext_ln1495_46_fu_1390_p1 = tmp_144_fu_1382_p3;

assign zext_ln1495_47_fu_1444_p1 = tmp_147_fu_1436_p3;

assign zext_ln1495_48_fu_1498_p1 = tmp_150_fu_1490_p3;

assign zext_ln1495_49_fu_1552_p1 = tmp_153_fu_1544_p3;

assign zext_ln1495_50_fu_1606_p1 = tmp_156_fu_1598_p3;

assign zext_ln1495_51_fu_1660_p1 = tmp_159_fu_1652_p3;

assign zext_ln1495_52_fu_1714_p1 = tmp_162_fu_1706_p3;

assign zext_ln1495_53_fu_1768_p1 = tmp_165_fu_1760_p3;

assign zext_ln1495_54_fu_1822_p1 = tmp_168_fu_1814_p3;

assign zext_ln1495_55_fu_1876_p1 = tmp_171_fu_1868_p3;

assign zext_ln1495_56_fu_1930_p1 = tmp_174_fu_1922_p3;

assign zext_ln1495_57_fu_1984_p1 = tmp_177_fu_1976_p3;

assign zext_ln1495_58_fu_2038_p1 = tmp_180_fu_2030_p3;

assign zext_ln1495_59_fu_2092_p1 = tmp_183_fu_2084_p3;

assign zext_ln1495_60_fu_2146_p1 = tmp_186_fu_2138_p3;

assign zext_ln1495_61_fu_2200_p1 = tmp_189_fu_2192_p3;

assign zext_ln1495_62_fu_2254_p1 = tmp_192_fu_2246_p3;

assign zext_ln1495_63_fu_2308_p1 = tmp_195_fu_2300_p3;

assign zext_ln1495_64_fu_2362_p1 = tmp_198_fu_2354_p3;

assign zext_ln1495_65_fu_2416_p1 = tmp_201_fu_2408_p3;

assign zext_ln1495_66_fu_2470_p1 = tmp_204_fu_2462_p3;

assign zext_ln1495_67_fu_2524_p1 = tmp_207_fu_2516_p3;

assign zext_ln1495_68_fu_2578_p1 = tmp_210_fu_2570_p3;

assign zext_ln1495_69_fu_2632_p1 = tmp_213_fu_2624_p3;

assign zext_ln1495_70_fu_2686_p1 = tmp_216_fu_2678_p3;

assign zext_ln1495_71_fu_2740_p1 = tmp_219_fu_2732_p3;

assign zext_ln1495_72_fu_2794_p1 = tmp_222_fu_2786_p3;

assign zext_ln1495_73_fu_2848_p1 = tmp_225_fu_2840_p3;

assign zext_ln1495_74_fu_2902_p1 = tmp_228_fu_2894_p3;

assign zext_ln1495_75_fu_2956_p1 = tmp_231_fu_2948_p3;

assign zext_ln1495_76_fu_3010_p1 = tmp_234_fu_3002_p3;

assign zext_ln1495_77_fu_3064_p1 = tmp_237_fu_3056_p3;

assign zext_ln1495_78_fu_3118_p1 = tmp_240_fu_3110_p3;

assign zext_ln1495_79_fu_3172_p1 = tmp_243_fu_3164_p3;

assign zext_ln1495_80_fu_3226_p1 = tmp_246_fu_3218_p3;

assign zext_ln1495_81_fu_3280_p1 = tmp_249_fu_3272_p3;

assign zext_ln1495_82_fu_3334_p1 = tmp_252_fu_3326_p3;

assign zext_ln1495_83_fu_3388_p1 = tmp_255_fu_3380_p3;

assign zext_ln1495_84_fu_3442_p1 = tmp_258_fu_3434_p3;

assign zext_ln1495_85_fu_3496_p1 = tmp_261_fu_3488_p3;

assign zext_ln1495_86_fu_3550_p1 = tmp_264_fu_3542_p3;

assign zext_ln1495_87_fu_3604_p1 = tmp_267_fu_3596_p3;

assign zext_ln1495_88_fu_3658_p1 = tmp_270_fu_3650_p3;

assign zext_ln1495_89_fu_3712_p1 = tmp_273_fu_3704_p3;

assign zext_ln1495_90_fu_3766_p1 = tmp_276_fu_3758_p3;

assign zext_ln1495_91_fu_3820_p1 = tmp_279_fu_3812_p3;

assign zext_ln1495_92_fu_3874_p1 = tmp_282_fu_3866_p3;

assign zext_ln1495_93_fu_3928_p1 = tmp_285_fu_3920_p3;

assign zext_ln1495_94_fu_3982_p1 = tmp_288_fu_3974_p3;

assign zext_ln1495_fu_580_p1 = tmp_99_fu_572_p3;

endmodule //relu_max_ap_fixed_ap_fixed_1_relu1_config5_s
// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and OpenCL
// Version: 2019.2
// Copyright (C) 1986-2019 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module relu_max_ap_fixed_ap_fixed_1_relu1_config9_s (
        ap_ready,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31
);


output   ap_ready;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;

wire   [0:0] tmp_2_fu_302_p3;
wire   [0:0] xor_ln1495_fu_310_p2;
wire   [10:0] tmp_3_fu_316_p3;
wire   [0:0] tmp_1_fu_288_p3;
wire   [0:0] icmp_ln1494_fu_296_p2;
wire   [0:0] or_ln1495_fu_328_p2;
wire   [15:0] zext_ln1495_fu_324_p1;
wire   [0:0] tmp_5_fu_356_p3;
wire   [0:0] xor_ln1495_1_fu_364_p2;
wire   [10:0] tmp_6_fu_370_p3;
wire   [0:0] tmp_4_fu_342_p3;
wire   [0:0] icmp_ln1494_1_fu_350_p2;
wire   [0:0] or_ln1495_1_fu_382_p2;
wire   [15:0] zext_ln1495_1_fu_378_p1;
wire   [0:0] tmp_8_fu_410_p3;
wire   [0:0] xor_ln1495_2_fu_418_p2;
wire   [10:0] tmp_9_fu_424_p3;
wire   [0:0] tmp_7_fu_396_p3;
wire   [0:0] icmp_ln1494_2_fu_404_p2;
wire   [0:0] or_ln1495_2_fu_436_p2;
wire   [15:0] zext_ln1495_2_fu_432_p1;
wire   [0:0] tmp_11_fu_464_p3;
wire   [0:0] xor_ln1495_3_fu_472_p2;
wire   [10:0] tmp_12_fu_478_p3;
wire   [0:0] tmp_10_fu_450_p3;
wire   [0:0] icmp_ln1494_3_fu_458_p2;
wire   [0:0] or_ln1495_3_fu_490_p2;
wire   [15:0] zext_ln1495_3_fu_486_p1;
wire   [0:0] tmp_14_fu_518_p3;
wire   [0:0] xor_ln1495_4_fu_526_p2;
wire   [10:0] tmp_15_fu_532_p3;
wire   [0:0] tmp_13_fu_504_p3;
wire   [0:0] icmp_ln1494_4_fu_512_p2;
wire   [0:0] or_ln1495_4_fu_544_p2;
wire   [15:0] zext_ln1495_4_fu_540_p1;
wire   [0:0] tmp_17_fu_572_p3;
wire   [0:0] xor_ln1495_5_fu_580_p2;
wire   [10:0] tmp_18_fu_586_p3;
wire   [0:0] tmp_16_fu_558_p3;
wire   [0:0] icmp_ln1494_5_fu_566_p2;
wire   [0:0] or_ln1495_5_fu_598_p2;
wire   [15:0] zext_ln1495_5_fu_594_p1;
wire   [0:0] tmp_20_fu_626_p3;
wire   [0:0] xor_ln1495_6_fu_634_p2;
wire   [10:0] tmp_21_fu_640_p3;
wire   [0:0] tmp_19_fu_612_p3;
wire   [0:0] icmp_ln1494_6_fu_620_p2;
wire   [0:0] or_ln1495_6_fu_652_p2;
wire   [15:0] zext_ln1495_6_fu_648_p1;
wire   [0:0] tmp_23_fu_680_p3;
wire   [0:0] xor_ln1495_7_fu_688_p2;
wire   [10:0] tmp_24_fu_694_p3;
wire   [0:0] tmp_22_fu_666_p3;
wire   [0:0] icmp_ln1494_7_fu_674_p2;
wire   [0:0] or_ln1495_7_fu_706_p2;
wire   [15:0] zext_ln1495_7_fu_702_p1;
wire   [0:0] tmp_26_fu_734_p3;
wire   [0:0] xor_ln1495_8_fu_742_p2;
wire   [10:0] tmp_27_fu_748_p3;
wire   [0:0] tmp_25_fu_720_p3;
wire   [0:0] icmp_ln1494_8_fu_728_p2;
wire   [0:0] or_ln1495_8_fu_760_p2;
wire   [15:0] zext_ln1495_8_fu_756_p1;
wire   [0:0] tmp_29_fu_788_p3;
wire   [0:0] xor_ln1495_9_fu_796_p2;
wire   [10:0] tmp_30_fu_802_p3;
wire   [0:0] tmp_28_fu_774_p3;
wire   [0:0] icmp_ln1494_9_fu_782_p2;
wire   [0:0] or_ln1495_9_fu_814_p2;
wire   [15:0] zext_ln1495_9_fu_810_p1;
wire   [0:0] tmp_32_fu_842_p3;
wire   [0:0] xor_ln1495_10_fu_850_p2;
wire   [10:0] tmp_33_fu_856_p3;
wire   [0:0] tmp_31_fu_828_p3;
wire   [0:0] icmp_ln1494_10_fu_836_p2;
wire   [0:0] or_ln1495_10_fu_868_p2;
wire   [15:0] zext_ln1495_10_fu_864_p1;
wire   [0:0] tmp_35_fu_896_p3;
wire   [0:0] xor_ln1495_11_fu_904_p2;
wire   [10:0] tmp_36_fu_910_p3;
wire   [0:0] tmp_34_fu_882_p3;
wire   [0:0] icmp_ln1494_11_fu_890_p2;
wire   [0:0] or_ln1495_11_fu_922_p2;
wire   [15:0] zext_ln1495_11_fu_918_p1;
wire   [0:0] tmp_38_fu_950_p3;
wire   [0:0] xor_ln1495_12_fu_958_p2;
wire   [10:0] tmp_39_fu_964_p3;
wire   [0:0] tmp_37_fu_936_p3;
wire   [0:0] icmp_ln1494_12_fu_944_p2;
wire   [0:0] or_ln1495_12_fu_976_p2;
wire   [15:0] zext_ln1495_12_fu_972_p1;
wire   [0:0] tmp_41_fu_1004_p3;
wire   [0:0] xor_ln1495_13_fu_1012_p2;
wire   [10:0] tmp_42_fu_1018_p3;
wire   [0:0] tmp_40_fu_990_p3;
wire   [0:0] icmp_ln1494_13_fu_998_p2;
wire   [0:0] or_ln1495_13_fu_1030_p2;
wire   [15:0] zext_ln1495_13_fu_1026_p1;
wire   [0:0] tmp_44_fu_1058_p3;
wire   [0:0] xor_ln1495_14_fu_1066_p2;
wire   [10:0] tmp_45_fu_1072_p3;
wire   [0:0] tmp_43_fu_1044_p3;
wire   [0:0] icmp_ln1494_14_fu_1052_p2;
wire   [0:0] or_ln1495_14_fu_1084_p2;
wire   [15:0] zext_ln1495_14_fu_1080_p1;
wire   [0:0] tmp_47_fu_1112_p3;
wire   [0:0] xor_ln1495_15_fu_1120_p2;
wire   [10:0] tmp_48_fu_1126_p3;
wire   [0:0] tmp_46_fu_1098_p3;
wire   [0:0] icmp_ln1494_15_fu_1106_p2;
wire   [0:0] or_ln1495_15_fu_1138_p2;
wire   [15:0] zext_ln1495_15_fu_1134_p1;
wire   [0:0] tmp_50_fu_1166_p3;
wire   [0:0] xor_ln1495_16_fu_1174_p2;
wire   [10:0] tmp_51_fu_1180_p3;
wire   [0:0] tmp_49_fu_1152_p3;
wire   [0:0] icmp_ln1494_16_fu_1160_p2;
wire   [0:0] or_ln1495_16_fu_1192_p2;
wire   [15:0] zext_ln1495_16_fu_1188_p1;
wire   [0:0] tmp_53_fu_1220_p3;
wire   [0:0] xor_ln1495_17_fu_1228_p2;
wire   [10:0] tmp_54_fu_1234_p3;
wire   [0:0] tmp_52_fu_1206_p3;
wire   [0:0] icmp_ln1494_17_fu_1214_p2;
wire   [0:0] or_ln1495_17_fu_1246_p2;
wire   [15:0] zext_ln1495_17_fu_1242_p1;
wire   [0:0] tmp_56_fu_1274_p3;
wire   [0:0] xor_ln1495_18_fu_1282_p2;
wire   [10:0] tmp_57_fu_1288_p3;
wire   [0:0] tmp_55_fu_1260_p3;
wire   [0:0] icmp_ln1494_18_fu_1268_p2;
wire   [0:0] or_ln1495_18_fu_1300_p2;
wire   [15:0] zext_ln1495_18_fu_1296_p1;
wire   [0:0] tmp_59_fu_1328_p3;
wire   [0:0] xor_ln1495_19_fu_1336_p2;
wire   [10:0] tmp_60_fu_1342_p3;
wire   [0:0] tmp_58_fu_1314_p3;
wire   [0:0] icmp_ln1494_19_fu_1322_p2;
wire   [0:0] or_ln1495_19_fu_1354_p2;
wire   [15:0] zext_ln1495_19_fu_1350_p1;
wire   [0:0] tmp_62_fu_1382_p3;
wire   [0:0] xor_ln1495_20_fu_1390_p2;
wire   [10:0] tmp_63_fu_1396_p3;
wire   [0:0] tmp_61_fu_1368_p3;
wire   [0:0] icmp_ln1494_20_fu_1376_p2;
wire   [0:0] or_ln1495_20_fu_1408_p2;
wire   [15:0] zext_ln1495_20_fu_1404_p1;
wire   [0:0] tmp_65_fu_1436_p3;
wire   [0:0] xor_ln1495_21_fu_1444_p2;
wire   [10:0] tmp_66_fu_1450_p3;
wire   [0:0] tmp_64_fu_1422_p3;
wire   [0:0] icmp_ln1494_21_fu_1430_p2;
wire   [0:0] or_ln1495_21_fu_1462_p2;
wire   [15:0] zext_ln1495_21_fu_1458_p1;
wire   [0:0] tmp_68_fu_1490_p3;
wire   [0:0] xor_ln1495_22_fu_1498_p2;
wire   [10:0] tmp_69_fu_1504_p3;
wire   [0:0] tmp_67_fu_1476_p3;
wire   [0:0] icmp_ln1494_22_fu_1484_p2;
wire   [0:0] or_ln1495_22_fu_1516_p2;
wire   [15:0] zext_ln1495_22_fu_1512_p1;
wire   [0:0] tmp_71_fu_1544_p3;
wire   [0:0] xor_ln1495_23_fu_1552_p2;
wire   [10:0] tmp_72_fu_1558_p3;
wire   [0:0] tmp_70_fu_1530_p3;
wire   [0:0] icmp_ln1494_23_fu_1538_p2;
wire   [0:0] or_ln1495_23_fu_1570_p2;
wire   [15:0] zext_ln1495_23_fu_1566_p1;
wire   [0:0] tmp_74_fu_1598_p3;
wire   [0:0] xor_ln1495_24_fu_1606_p2;
wire   [10:0] tmp_75_fu_1612_p3;
wire   [0:0] tmp_73_fu_1584_p3;
wire   [0:0] icmp_ln1494_24_fu_1592_p2;
wire   [0:0] or_ln1495_24_fu_1624_p2;
wire   [15:0] zext_ln1495_24_fu_1620_p1;
wire   [0:0] tmp_77_fu_1652_p3;
wire   [0:0] xor_ln1495_25_fu_1660_p2;
wire   [10:0] tmp_78_fu_1666_p3;
wire   [0:0] tmp_76_fu_1638_p3;
wire   [0:0] icmp_ln1494_25_fu_1646_p2;
wire   [0:0] or_ln1495_25_fu_1678_p2;
wire   [15:0] zext_ln1495_25_fu_1674_p1;
wire   [0:0] tmp_80_fu_1706_p3;
wire   [0:0] xor_ln1495_26_fu_1714_p2;
wire   [10:0] tmp_81_fu_1720_p3;
wire   [0:0] tmp_79_fu_1692_p3;
wire   [0:0] icmp_ln1494_26_fu_1700_p2;
wire   [0:0] or_ln1495_26_fu_1732_p2;
wire   [15:0] zext_ln1495_26_fu_1728_p1;
wire   [0:0] tmp_83_fu_1760_p3;
wire   [0:0] xor_ln1495_27_fu_1768_p2;
wire   [10:0] tmp_84_fu_1774_p3;
wire   [0:0] tmp_82_fu_1746_p3;
wire   [0:0] icmp_ln1494_27_fu_1754_p2;
wire   [0:0] or_ln1495_27_fu_1786_p2;
wire   [15:0] zext_ln1495_27_fu_1782_p1;
wire   [0:0] tmp_86_fu_1814_p3;
wire   [0:0] xor_ln1495_28_fu_1822_p2;
wire   [10:0] tmp_87_fu_1828_p3;
wire   [0:0] tmp_85_fu_1800_p3;
wire   [0:0] icmp_ln1494_28_fu_1808_p2;
wire   [0:0] or_ln1495_28_fu_1840_p2;
wire   [15:0] zext_ln1495_28_fu_1836_p1;
wire   [0:0] tmp_89_fu_1868_p3;
wire   [0:0] xor_ln1495_29_fu_1876_p2;
wire   [10:0] tmp_90_fu_1882_p3;
wire   [0:0] tmp_88_fu_1854_p3;
wire   [0:0] icmp_ln1494_29_fu_1862_p2;
wire   [0:0] or_ln1495_29_fu_1894_p2;
wire   [15:0] zext_ln1495_29_fu_1890_p1;
wire   [0:0] tmp_92_fu_1922_p3;
wire   [0:0] xor_ln1495_30_fu_1930_p2;
wire   [10:0] tmp_93_fu_1936_p3;
wire   [0:0] tmp_91_fu_1908_p3;
wire   [0:0] icmp_ln1494_30_fu_1916_p2;
wire   [0:0] or_ln1495_30_fu_1948_p2;
wire   [15:0] zext_ln1495_30_fu_1944_p1;
wire   [0:0] tmp_95_fu_1976_p3;
wire   [0:0] xor_ln1495_31_fu_1984_p2;
wire   [10:0] tmp_96_fu_1990_p3;
wire   [0:0] tmp_94_fu_1962_p3;
wire   [0:0] icmp_ln1494_31_fu_1970_p2;
wire   [0:0] or_ln1495_31_fu_2002_p2;
wire   [15:0] zext_ln1495_31_fu_1998_p1;
wire   [15:0] select_ln1495_fu_334_p3;
wire   [15:0] select_ln1495_1_fu_388_p3;
wire   [15:0] select_ln1495_2_fu_442_p3;
wire   [15:0] select_ln1495_3_fu_496_p3;
wire   [15:0] select_ln1495_4_fu_550_p3;
wire   [15:0] select_ln1495_5_fu_604_p3;
wire   [15:0] select_ln1495_6_fu_658_p3;
wire   [15:0] select_ln1495_7_fu_712_p3;
wire   [15:0] select_ln1495_8_fu_766_p3;
wire   [15:0] select_ln1495_9_fu_820_p3;
wire   [15:0] select_ln1495_10_fu_874_p3;
wire   [15:0] select_ln1495_11_fu_928_p3;
wire   [15:0] select_ln1495_12_fu_982_p3;
wire   [15:0] select_ln1495_13_fu_1036_p3;
wire   [15:0] select_ln1495_14_fu_1090_p3;
wire   [15:0] select_ln1495_15_fu_1144_p3;
wire   [15:0] select_ln1495_16_fu_1198_p3;
wire   [15:0] select_ln1495_17_fu_1252_p3;
wire   [15:0] select_ln1495_18_fu_1306_p3;
wire   [15:0] select_ln1495_19_fu_1360_p3;
wire   [15:0] select_ln1495_20_fu_1414_p3;
wire   [15:0] select_ln1495_21_fu_1468_p3;
wire   [15:0] select_ln1495_22_fu_1522_p3;
wire   [15:0] select_ln1495_23_fu_1576_p3;
wire   [15:0] select_ln1495_24_fu_1630_p3;
wire   [15:0] select_ln1495_25_fu_1684_p3;
wire   [15:0] select_ln1495_26_fu_1738_p3;
wire   [15:0] select_ln1495_27_fu_1792_p3;
wire   [15:0] select_ln1495_28_fu_1846_p3;
wire   [15:0] select_ln1495_29_fu_1900_p3;
wire   [15:0] select_ln1495_30_fu_1954_p3;
wire   [15:0] select_ln1495_31_fu_2008_p3;

assign ap_ready = 1'b1;

assign ap_return_0 = select_ln1495_fu_334_p3;

assign ap_return_1 = select_ln1495_1_fu_388_p3;

assign ap_return_10 = select_ln1495_10_fu_874_p3;

assign ap_return_11 = select_ln1495_11_fu_928_p3;

assign ap_return_12 = select_ln1495_12_fu_982_p3;

assign ap_return_13 = select_ln1495_13_fu_1036_p3;

assign ap_return_14 = select_ln1495_14_fu_1090_p3;

assign ap_return_15 = select_ln1495_15_fu_1144_p3;

assign ap_return_16 = select_ln1495_16_fu_1198_p3;

assign ap_return_17 = select_ln1495_17_fu_1252_p3;

assign ap_return_18 = select_ln1495_18_fu_1306_p3;

assign ap_return_19 = select_ln1495_19_fu_1360_p3;

assign ap_return_2 = select_ln1495_2_fu_442_p3;

assign ap_return_20 = select_ln1495_20_fu_1414_p3;

assign ap_return_21 = select_ln1495_21_fu_1468_p3;

assign ap_return_22 = select_ln1495_22_fu_1522_p3;

assign ap_return_23 = select_ln1495_23_fu_1576_p3;

assign ap_return_24 = select_ln1495_24_fu_1630_p3;

assign ap_return_25 = select_ln1495_25_fu_1684_p3;

assign ap_return_26 = select_ln1495_26_fu_1738_p3;

assign ap_return_27 = select_ln1495_27_fu_1792_p3;

assign ap_return_28 = select_ln1495_28_fu_1846_p3;

assign ap_return_29 = select_ln1495_29_fu_1900_p3;

assign ap_return_3 = select_ln1495_3_fu_496_p3;

assign ap_return_30 = select_ln1495_30_fu_1954_p3;

assign ap_return_31 = select_ln1495_31_fu_2008_p3;

assign ap_return_4 = select_ln1495_4_fu_550_p3;

assign ap_return_5 = select_ln1495_5_fu_604_p3;

assign ap_return_6 = select_ln1495_6_fu_658_p3;

assign ap_return_7 = select_ln1495_7_fu_712_p3;

assign ap_return_8 = select_ln1495_8_fu_766_p3;

assign ap_return_9 = select_ln1495_9_fu_820_p3;

assign icmp_ln1494_10_fu_836_p2 = (((data_10_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_11_fu_890_p2 = (((data_11_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_12_fu_944_p2 = (((data_12_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_13_fu_998_p2 = (((data_13_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_14_fu_1052_p2 = (((data_14_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_15_fu_1106_p2 = (((data_15_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_16_fu_1160_p2 = (((data_16_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_17_fu_1214_p2 = (((data_17_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_18_fu_1268_p2 = (((data_18_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_19_fu_1322_p2 = (((data_19_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_1_fu_350_p2 = (((data_1_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_20_fu_1376_p2 = (((data_20_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_21_fu_1430_p2 = (((data_21_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_22_fu_1484_p2 = (((data_22_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_23_fu_1538_p2 = (((data_23_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_24_fu_1592_p2 = (((data_24_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_25_fu_1646_p2 = (((data_25_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_26_fu_1700_p2 = (((data_26_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_27_fu_1754_p2 = (((data_27_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_28_fu_1808_p2 = (((data_28_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_29_fu_1862_p2 = (((data_29_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_2_fu_404_p2 = (((data_2_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_30_fu_1916_p2 = (((data_30_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_31_fu_1970_p2 = (((data_31_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_3_fu_458_p2 = (((data_3_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_4_fu_512_p2 = (((data_4_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_5_fu_566_p2 = (((data_5_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_6_fu_620_p2 = (((data_6_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_7_fu_674_p2 = (((data_7_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_8_fu_728_p2 = (((data_8_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_9_fu_782_p2 = (((data_9_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_fu_296_p2 = (((data_0_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign or_ln1495_10_fu_868_p2 = (tmp_31_fu_828_p3 | icmp_ln1494_10_fu_836_p2);

assign or_ln1495_11_fu_922_p2 = (tmp_34_fu_882_p3 | icmp_ln1494_11_fu_890_p2);

assign or_ln1495_12_fu_976_p2 = (tmp_37_fu_936_p3 | icmp_ln1494_12_fu_944_p2);

assign or_ln1495_13_fu_1030_p2 = (tmp_40_fu_990_p3 | icmp_ln1494_13_fu_998_p2);

assign or_ln1495_14_fu_1084_p2 = (tmp_43_fu_1044_p3 | icmp_ln1494_14_fu_1052_p2);

assign or_ln1495_15_fu_1138_p2 = (tmp_46_fu_1098_p3 | icmp_ln1494_15_fu_1106_p2);

assign or_ln1495_16_fu_1192_p2 = (tmp_49_fu_1152_p3 | icmp_ln1494_16_fu_1160_p2);

assign or_ln1495_17_fu_1246_p2 = (tmp_52_fu_1206_p3 | icmp_ln1494_17_fu_1214_p2);

assign or_ln1495_18_fu_1300_p2 = (tmp_55_fu_1260_p3 | icmp_ln1494_18_fu_1268_p2);

assign or_ln1495_19_fu_1354_p2 = (tmp_58_fu_1314_p3 | icmp_ln1494_19_fu_1322_p2);

assign or_ln1495_1_fu_382_p2 = (tmp_4_fu_342_p3 | icmp_ln1494_1_fu_350_p2);

assign or_ln1495_20_fu_1408_p2 = (tmp_61_fu_1368_p3 | icmp_ln1494_20_fu_1376_p2);

assign or_ln1495_21_fu_1462_p2 = (tmp_64_fu_1422_p3 | icmp_ln1494_21_fu_1430_p2);

assign or_ln1495_22_fu_1516_p2 = (tmp_67_fu_1476_p3 | icmp_ln1494_22_fu_1484_p2);

assign or_ln1495_23_fu_1570_p2 = (tmp_70_fu_1530_p3 | icmp_ln1494_23_fu_1538_p2);

assign or_ln1495_24_fu_1624_p2 = (tmp_73_fu_1584_p3 | icmp_ln1494_24_fu_1592_p2);

assign or_ln1495_25_fu_1678_p2 = (tmp_76_fu_1638_p3 | icmp_ln1494_25_fu_1646_p2);

assign or_ln1495_26_fu_1732_p2 = (tmp_79_fu_1692_p3 | icmp_ln1494_26_fu_1700_p2);

assign or_ln1495_27_fu_1786_p2 = (tmp_82_fu_1746_p3 | icmp_ln1494_27_fu_1754_p2);

assign or_ln1495_28_fu_1840_p2 = (tmp_85_fu_1800_p3 | icmp_ln1494_28_fu_1808_p2);

assign or_ln1495_29_fu_1894_p2 = (tmp_88_fu_1854_p3 | icmp_ln1494_29_fu_1862_p2);

assign or_ln1495_2_fu_436_p2 = (tmp_7_fu_396_p3 | icmp_ln1494_2_fu_404_p2);

assign or_ln1495_30_fu_1948_p2 = (tmp_91_fu_1908_p3 | icmp_ln1494_30_fu_1916_p2);

assign or_ln1495_31_fu_2002_p2 = (tmp_94_fu_1962_p3 | icmp_ln1494_31_fu_1970_p2);

assign or_ln1495_3_fu_490_p2 = (tmp_10_fu_450_p3 | icmp_ln1494_3_fu_458_p2);

assign or_ln1495_4_fu_544_p2 = (tmp_13_fu_504_p3 | icmp_ln1494_4_fu_512_p2);

assign or_ln1495_5_fu_598_p2 = (tmp_16_fu_558_p3 | icmp_ln1494_5_fu_566_p2);

assign or_ln1495_6_fu_652_p2 = (tmp_19_fu_612_p3 | icmp_ln1494_6_fu_620_p2);

assign or_ln1495_7_fu_706_p2 = (tmp_22_fu_666_p3 | icmp_ln1494_7_fu_674_p2);

assign or_ln1495_8_fu_760_p2 = (tmp_25_fu_720_p3 | icmp_ln1494_8_fu_728_p2);

assign or_ln1495_9_fu_814_p2 = (tmp_28_fu_774_p3 | icmp_ln1494_9_fu_782_p2);

assign or_ln1495_fu_328_p2 = (tmp_1_fu_288_p3 | icmp_ln1494_fu_296_p2);

assign select_ln1495_10_fu_874_p3 = ((or_ln1495_10_fu_868_p2[0:0] == 1'b1) ? zext_ln1495_10_fu_864_p1 : data_10_V_read);

assign select_ln1495_11_fu_928_p3 = ((or_ln1495_11_fu_922_p2[0:0] == 1'b1) ? zext_ln1495_11_fu_918_p1 : data_11_V_read);

assign select_ln1495_12_fu_982_p3 = ((or_ln1495_12_fu_976_p2[0:0] == 1'b1) ? zext_ln1495_12_fu_972_p1 : data_12_V_read);

assign select_ln1495_13_fu_1036_p3 = ((or_ln1495_13_fu_1030_p2[0:0] == 1'b1) ? zext_ln1495_13_fu_1026_p1 : data_13_V_read);

assign select_ln1495_14_fu_1090_p3 = ((or_ln1495_14_fu_1084_p2[0:0] == 1'b1) ? zext_ln1495_14_fu_1080_p1 : data_14_V_read);

assign select_ln1495_15_fu_1144_p3 = ((or_ln1495_15_fu_1138_p2[0:0] == 1'b1) ? zext_ln1495_15_fu_1134_p1 : data_15_V_read);

assign select_ln1495_16_fu_1198_p3 = ((or_ln1495_16_fu_1192_p2[0:0] == 1'b1) ? zext_ln1495_16_fu_1188_p1 : data_16_V_read);

assign select_ln1495_17_fu_1252_p3 = ((or_ln1495_17_fu_1246_p2[0:0] == 1'b1) ? zext_ln1495_17_fu_1242_p1 : data_17_V_read);

assign select_ln1495_18_fu_1306_p3 = ((or_ln1495_18_fu_1300_p2[0:0] == 1'b1) ? zext_ln1495_18_fu_1296_p1 : data_18_V_read);

assign select_ln1495_19_fu_1360_p3 = ((or_ln1495_19_fu_1354_p2[0:0] == 1'b1) ? zext_ln1495_19_fu_1350_p1 : data_19_V_read);

assign select_ln1495_1_fu_388_p3 = ((or_ln1495_1_fu_382_p2[0:0] == 1'b1) ? zext_ln1495_1_fu_378_p1 : data_1_V_read);

assign select_ln1495_20_fu_1414_p3 = ((or_ln1495_20_fu_1408_p2[0:0] == 1'b1) ? zext_ln1495_20_fu_1404_p1 : data_20_V_read);

assign select_ln1495_21_fu_1468_p3 = ((or_ln1495_21_fu_1462_p2[0:0] == 1'b1) ? zext_ln1495_21_fu_1458_p1 : data_21_V_read);

assign select_ln1495_22_fu_1522_p3 = ((or_ln1495_22_fu_1516_p2[0:0] == 1'b1) ? zext_ln1495_22_fu_1512_p1 : data_22_V_read);

assign select_ln1495_23_fu_1576_p3 = ((or_ln1495_23_fu_1570_p2[0:0] == 1'b1) ? zext_ln1495_23_fu_1566_p1 : data_23_V_read);

assign select_ln1495_24_fu_1630_p3 = ((or_ln1495_24_fu_1624_p2[0:0] == 1'b1) ? zext_ln1495_24_fu_1620_p1 : data_24_V_read);

assign select_ln1495_25_fu_1684_p3 = ((or_ln1495_25_fu_1678_p2[0:0] == 1'b1) ? zext_ln1495_25_fu_1674_p1 : data_25_V_read);

assign select_ln1495_26_fu_1738_p3 = ((or_ln1495_26_fu_1732_p2[0:0] == 1'b1) ? zext_ln1495_26_fu_1728_p1 : data_26_V_read);

assign select_ln1495_27_fu_1792_p3 = ((or_ln1495_27_fu_1786_p2[0:0] == 1'b1) ? zext_ln1495_27_fu_1782_p1 : data_27_V_read);

assign select_ln1495_28_fu_1846_p3 = ((or_ln1495_28_fu_1840_p2[0:0] == 1'b1) ? zext_ln1495_28_fu_1836_p1 : data_28_V_read);

assign select_ln1495_29_fu_1900_p3 = ((or_ln1495_29_fu_1894_p2[0:0] == 1'b1) ? zext_ln1495_29_fu_1890_p1 : data_29_V_read);

assign select_ln1495_2_fu_442_p3 = ((or_ln1495_2_fu_436_p2[0:0] == 1'b1) ? zext_ln1495_2_fu_432_p1 : data_2_V_read);

assign select_ln1495_30_fu_1954_p3 = ((or_ln1495_30_fu_1948_p2[0:0] == 1'b1) ? zext_ln1495_30_fu_1944_p1 : data_30_V_read);

assign select_ln1495_31_fu_2008_p3 = ((or_ln1495_31_fu_2002_p2[0:0] == 1'b1) ? zext_ln1495_31_fu_1998_p1 : data_31_V_read);

assign select_ln1495_3_fu_496_p3 = ((or_ln1495_3_fu_490_p2[0:0] == 1'b1) ? zext_ln1495_3_fu_486_p1 : data_3_V_read);

assign select_ln1495_4_fu_550_p3 = ((or_ln1495_4_fu_544_p2[0:0] == 1'b1) ? zext_ln1495_4_fu_540_p1 : data_4_V_read);

assign select_ln1495_5_fu_604_p3 = ((or_ln1495_5_fu_598_p2[0:0] == 1'b1) ? zext_ln1495_5_fu_594_p1 : data_5_V_read);

assign select_ln1495_6_fu_658_p3 = ((or_ln1495_6_fu_652_p2[0:0] == 1'b1) ? zext_ln1495_6_fu_648_p1 : data_6_V_read);

assign select_ln1495_7_fu_712_p3 = ((or_ln1495_7_fu_706_p2[0:0] == 1'b1) ? zext_ln1495_7_fu_702_p1 : data_7_V_read);

assign select_ln1495_8_fu_766_p3 = ((or_ln1495_8_fu_760_p2[0:0] == 1'b1) ? zext_ln1495_8_fu_756_p1 : data_8_V_read);

assign select_ln1495_9_fu_820_p3 = ((or_ln1495_9_fu_814_p2[0:0] == 1'b1) ? zext_ln1495_9_fu_810_p1 : data_9_V_read);

assign select_ln1495_fu_334_p3 = ((or_ln1495_fu_328_p2[0:0] == 1'b1) ? zext_ln1495_fu_324_p1 : data_0_V_read);

assign tmp_10_fu_450_p3 = data_3_V_read[32'd15];

assign tmp_11_fu_464_p3 = data_3_V_read[32'd15];

assign tmp_12_fu_478_p3 = {{xor_ln1495_3_fu_472_p2}, {10'd0}};

assign tmp_13_fu_504_p3 = data_4_V_read[32'd15];

assign tmp_14_fu_518_p3 = data_4_V_read[32'd15];

assign tmp_15_fu_532_p3 = {{xor_ln1495_4_fu_526_p2}, {10'd0}};

assign tmp_16_fu_558_p3 = data_5_V_read[32'd15];

assign tmp_17_fu_572_p3 = data_5_V_read[32'd15];

assign tmp_18_fu_586_p3 = {{xor_ln1495_5_fu_580_p2}, {10'd0}};

assign tmp_19_fu_612_p3 = data_6_V_read[32'd15];

assign tmp_1_fu_288_p3 = data_0_V_read[32'd15];

assign tmp_20_fu_626_p3 = data_6_V_read[32'd15];

assign tmp_21_fu_640_p3 = {{xor_ln1495_6_fu_634_p2}, {10'd0}};

assign tmp_22_fu_666_p3 = data_7_V_read[32'd15];

assign tmp_23_fu_680_p3 = data_7_V_read[32'd15];

assign tmp_24_fu_694_p3 = {{xor_ln1495_7_fu_688_p2}, {10'd0}};

assign tmp_25_fu_720_p3 = data_8_V_read[32'd15];

assign tmp_26_fu_734_p3 = data_8_V_read[32'd15];

assign tmp_27_fu_748_p3 = {{xor_ln1495_8_fu_742_p2}, {10'd0}};

assign tmp_28_fu_774_p3 = data_9_V_read[32'd15];

assign tmp_29_fu_788_p3 = data_9_V_read[32'd15];

assign tmp_2_fu_302_p3 = data_0_V_read[32'd15];

assign tmp_30_fu_802_p3 = {{xor_ln1495_9_fu_796_p2}, {10'd0}};

assign tmp_31_fu_828_p3 = data_10_V_read[32'd15];

assign tmp_32_fu_842_p3 = data_10_V_read[32'd15];

assign tmp_33_fu_856_p3 = {{xor_ln1495_10_fu_850_p2}, {10'd0}};

assign tmp_34_fu_882_p3 = data_11_V_read[32'd15];

assign tmp_35_fu_896_p3 = data_11_V_read[32'd15];

assign tmp_36_fu_910_p3 = {{xor_ln1495_11_fu_904_p2}, {10'd0}};

assign tmp_37_fu_936_p3 = data_12_V_read[32'd15];

assign tmp_38_fu_950_p3 = data_12_V_read[32'd15];

assign tmp_39_fu_964_p3 = {{xor_ln1495_12_fu_958_p2}, {10'd0}};

assign tmp_3_fu_316_p3 = {{xor_ln1495_fu_310_p2}, {10'd0}};

assign tmp_40_fu_990_p3 = data_13_V_read[32'd15];

assign tmp_41_fu_1004_p3 = data_13_V_read[32'd15];

assign tmp_42_fu_1018_p3 = {{xor_ln1495_13_fu_1012_p2}, {10'd0}};

assign tmp_43_fu_1044_p3 = data_14_V_read[32'd15];

assign tmp_44_fu_1058_p3 = data_14_V_read[32'd15];

assign tmp_45_fu_1072_p3 = {{xor_ln1495_14_fu_1066_p2}, {10'd0}};

assign tmp_46_fu_1098_p3 = data_15_V_read[32'd15];

assign tmp_47_fu_1112_p3 = data_15_V_read[32'd15];

assign tmp_48_fu_1126_p3 = {{xor_ln1495_15_fu_1120_p2}, {10'd0}};

assign tmp_49_fu_1152_p3 = data_16_V_read[32'd15];

assign tmp_4_fu_342_p3 = data_1_V_read[32'd15];

assign tmp_50_fu_1166_p3 = data_16_V_read[32'd15];

assign tmp_51_fu_1180_p3 = {{xor_ln1495_16_fu_1174_p2}, {10'd0}};

assign tmp_52_fu_1206_p3 = data_17_V_read[32'd15];

assign tmp_53_fu_1220_p3 = data_17_V_read[32'd15];

assign tmp_54_fu_1234_p3 = {{xor_ln1495_17_fu_1228_p2}, {10'd0}};

assign tmp_55_fu_1260_p3 = data_18_V_read[32'd15];

assign tmp_56_fu_1274_p3 = data_18_V_read[32'd15];

assign tmp_57_fu_1288_p3 = {{xor_ln1495_18_fu_1282_p2}, {10'd0}};

assign tmp_58_fu_1314_p3 = data_19_V_read[32'd15];

assign tmp_59_fu_1328_p3 = data_19_V_read[32'd15];

assign tmp_5_fu_356_p3 = data_1_V_read[32'd15];

assign tmp_60_fu_1342_p3 = {{xor_ln1495_19_fu_1336_p2}, {10'd0}};

assign tmp_61_fu_1368_p3 = data_20_V_read[32'd15];

assign tmp_62_fu_1382_p3 = data_20_V_read[32'd15];

assign tmp_63_fu_1396_p3 = {{xor_ln1495_20_fu_1390_p2}, {10'd0}};

assign tmp_64_fu_1422_p3 = data_21_V_read[32'd15];

assign tmp_65_fu_1436_p3 = data_21_V_read[32'd15];

assign tmp_66_fu_1450_p3 = {{xor_ln1495_21_fu_1444_p2}, {10'd0}};

assign tmp_67_fu_1476_p3 = data_22_V_read[32'd15];

assign tmp_68_fu_1490_p3 = data_22_V_read[32'd15];

assign tmp_69_fu_1504_p3 = {{xor_ln1495_22_fu_1498_p2}, {10'd0}};

assign tmp_6_fu_370_p3 = {{xor_ln1495_1_fu_364_p2}, {10'd0}};

assign tmp_70_fu_1530_p3 = data_23_V_read[32'd15];

assign tmp_71_fu_1544_p3 = data_23_V_read[32'd15];

assign tmp_72_fu_1558_p3 = {{xor_ln1495_23_fu_1552_p2}, {10'd0}};

assign tmp_73_fu_1584_p3 = data_24_V_read[32'd15];

assign tmp_74_fu_1598_p3 = data_24_V_read[32'd15];

assign tmp_75_fu_1612_p3 = {{xor_ln1495_24_fu_1606_p2}, {10'd0}};

assign tmp_76_fu_1638_p3 = data_25_V_read[32'd15];

assign tmp_77_fu_1652_p3 = data_25_V_read[32'd15];

assign tmp_78_fu_1666_p3 = {{xor_ln1495_25_fu_1660_p2}, {10'd0}};

assign tmp_79_fu_1692_p3 = data_26_V_read[32'd15];

assign tmp_7_fu_396_p3 = data_2_V_read[32'd15];

assign tmp_80_fu_1706_p3 = data_26_V_read[32'd15];

assign tmp_81_fu_1720_p3 = {{xor_ln1495_26_fu_1714_p2}, {10'd0}};

assign tmp_82_fu_1746_p3 = data_27_V_read[32'd15];

assign tmp_83_fu_1760_p3 = data_27_V_read[32'd15];

assign tmp_84_fu_1774_p3 = {{xor_ln1495_27_fu_1768_p2}, {10'd0}};

assign tmp_85_fu_1800_p3 = data_28_V_read[32'd15];

assign tmp_86_fu_1814_p3 = data_28_V_read[32'd15];

assign tmp_87_fu_1828_p3 = {{xor_ln1495_28_fu_1822_p2}, {10'd0}};

assign tmp_88_fu_1854_p3 = data_29_V_read[32'd15];

assign tmp_89_fu_1868_p3 = data_29_V_read[32'd15];

assign tmp_8_fu_410_p3 = data_2_V_read[32'd15];

assign tmp_90_fu_1882_p3 = {{xor_ln1495_29_fu_1876_p2}, {10'd0}};

assign tmp_91_fu_1908_p3 = data_30_V_read[32'd15];

assign tmp_92_fu_1922_p3 = data_30_V_read[32'd15];

assign tmp_93_fu_1936_p3 = {{xor_ln1495_30_fu_1930_p2}, {10'd0}};

assign tmp_94_fu_1962_p3 = data_31_V_read[32'd15];

assign tmp_95_fu_1976_p3 = data_31_V_read[32'd15];

assign tmp_96_fu_1990_p3 = {{xor_ln1495_31_fu_1984_p2}, {10'd0}};

assign tmp_9_fu_424_p3 = {{xor_ln1495_2_fu_418_p2}, {10'd0}};

assign xor_ln1495_10_fu_850_p2 = (tmp_32_fu_842_p3 ^ 1'd1);

assign xor_ln1495_11_fu_904_p2 = (tmp_35_fu_896_p3 ^ 1'd1);

assign xor_ln1495_12_fu_958_p2 = (tmp_38_fu_950_p3 ^ 1'd1);

assign xor_ln1495_13_fu_1012_p2 = (tmp_41_fu_1004_p3 ^ 1'd1);

assign xor_ln1495_14_fu_1066_p2 = (tmp_44_fu_1058_p3 ^ 1'd1);

assign xor_ln1495_15_fu_1120_p2 = (tmp_47_fu_1112_p3 ^ 1'd1);

assign xor_ln1495_16_fu_1174_p2 = (tmp_50_fu_1166_p3 ^ 1'd1);

assign xor_ln1495_17_fu_1228_p2 = (tmp_53_fu_1220_p3 ^ 1'd1);

assign xor_ln1495_18_fu_1282_p2 = (tmp_56_fu_1274_p3 ^ 1'd1);

assign xor_ln1495_19_fu_1336_p2 = (tmp_59_fu_1328_p3 ^ 1'd1);

assign xor_ln1495_1_fu_364_p2 = (tmp_5_fu_356_p3 ^ 1'd1);

assign xor_ln1495_20_fu_1390_p2 = (tmp_62_fu_1382_p3 ^ 1'd1);

assign xor_ln1495_21_fu_1444_p2 = (tmp_65_fu_1436_p3 ^ 1'd1);

assign xor_ln1495_22_fu_1498_p2 = (tmp_68_fu_1490_p3 ^ 1'd1);

assign xor_ln1495_23_fu_1552_p2 = (tmp_71_fu_1544_p3 ^ 1'd1);

assign xor_ln1495_24_fu_1606_p2 = (tmp_74_fu_1598_p3 ^ 1'd1);

assign xor_ln1495_25_fu_1660_p2 = (tmp_77_fu_1652_p3 ^ 1'd1);

assign xor_ln1495_26_fu_1714_p2 = (tmp_80_fu_1706_p3 ^ 1'd1);

assign xor_ln1495_27_fu_1768_p2 = (tmp_83_fu_1760_p3 ^ 1'd1);

assign xor_ln1495_28_fu_1822_p2 = (tmp_86_fu_1814_p3 ^ 1'd1);

assign xor_ln1495_29_fu_1876_p2 = (tmp_89_fu_1868_p3 ^ 1'd1);

assign xor_ln1495_2_fu_418_p2 = (tmp_8_fu_410_p3 ^ 1'd1);

assign xor_ln1495_30_fu_1930_p2 = (tmp_92_fu_1922_p3 ^ 1'd1);

assign xor_ln1495_31_fu_1984_p2 = (tmp_95_fu_1976_p3 ^ 1'd1);

assign xor_ln1495_3_fu_472_p2 = (tmp_11_fu_464_p3 ^ 1'd1);

assign xor_ln1495_4_fu_526_p2 = (tmp_14_fu_518_p3 ^ 1'd1);

assign xor_ln1495_5_fu_580_p2 = (tmp_17_fu_572_p3 ^ 1'd1);

assign xor_ln1495_6_fu_634_p2 = (tmp_20_fu_626_p3 ^ 1'd1);

assign xor_ln1495_7_fu_688_p2 = (tmp_23_fu_680_p3 ^ 1'd1);

assign xor_ln1495_8_fu_742_p2 = (tmp_26_fu_734_p3 ^ 1'd1);

assign xor_ln1495_9_fu_796_p2 = (tmp_29_fu_788_p3 ^ 1'd1);

assign xor_ln1495_fu_310_p2 = (tmp_2_fu_302_p3 ^ 1'd1);

assign zext_ln1495_10_fu_864_p1 = tmp_33_fu_856_p3;

assign zext_ln1495_11_fu_918_p1 = tmp_36_fu_910_p3;

assign zext_ln1495_12_fu_972_p1 = tmp_39_fu_964_p3;

assign zext_ln1495_13_fu_1026_p1 = tmp_42_fu_1018_p3;

assign zext_ln1495_14_fu_1080_p1 = tmp_45_fu_1072_p3;

assign zext_ln1495_15_fu_1134_p1 = tmp_48_fu_1126_p3;

assign zext_ln1495_16_fu_1188_p1 = tmp_51_fu_1180_p3;

assign zext_ln1495_17_fu_1242_p1 = tmp_54_fu_1234_p3;

assign zext_ln1495_18_fu_1296_p1 = tmp_57_fu_1288_p3;

assign zext_ln1495_19_fu_1350_p1 = tmp_60_fu_1342_p3;

assign zext_ln1495_1_fu_378_p1 = tmp_6_fu_370_p3;

assign zext_ln1495_20_fu_1404_p1 = tmp_63_fu_1396_p3;

assign zext_ln1495_21_fu_1458_p1 = tmp_66_fu_1450_p3;

assign zext_ln1495_22_fu_1512_p1 = tmp_69_fu_1504_p3;

assign zext_ln1495_23_fu_1566_p1 = tmp_72_fu_1558_p3;

assign zext_ln1495_24_fu_1620_p1 = tmp_75_fu_1612_p3;

assign zext_ln1495_25_fu_1674_p1 = tmp_78_fu_1666_p3;

assign zext_ln1495_26_fu_1728_p1 = tmp_81_fu_1720_p3;

assign zext_ln1495_27_fu_1782_p1 = tmp_84_fu_1774_p3;

assign zext_ln1495_28_fu_1836_p1 = tmp_87_fu_1828_p3;

assign zext_ln1495_29_fu_1890_p1 = tmp_90_fu_1882_p3;

assign zext_ln1495_2_fu_432_p1 = tmp_9_fu_424_p3;

assign zext_ln1495_30_fu_1944_p1 = tmp_93_fu_1936_p3;

assign zext_ln1495_31_fu_1998_p1 = tmp_96_fu_1990_p3;

assign zext_ln1495_3_fu_486_p1 = tmp_12_fu_478_p3;

assign zext_ln1495_4_fu_540_p1 = tmp_15_fu_532_p3;

assign zext_ln1495_5_fu_594_p1 = tmp_18_fu_586_p3;

assign zext_ln1495_6_fu_648_p1 = tmp_21_fu_640_p3;

assign zext_ln1495_7_fu_702_p1 = tmp_24_fu_694_p3;

assign zext_ln1495_8_fu_756_p1 = tmp_27_fu_748_p3;

assign zext_ln1495_9_fu_810_p1 = tmp_30_fu_802_p3;

assign zext_ln1495_fu_324_p1 = tmp_3_fu_316_p3;

endmodule //relu_max_ap_fixed_ap_fixed_1_relu1_config9_s
