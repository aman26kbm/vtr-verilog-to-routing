`define BRAM_DWIDTH 40
`define BRAM_AWIDTH 9
`define BRAM_DEPTH 512
`define COMPUTE_DWIDTH 4
`define NUM 10

module system(
  input clk,
  input reset,
  input start,
  output done,
  input external,
  input  [`BRAM_AWIDTH-1:0] bram_addr_ext,
  output [`BRAM_DWIDTH-1:0] bram_rdata_ext,
  input  [`BRAM_DWIDTH-1:0] bram_wdata_ext,
  input  bram_wren_ext,
  input [`BRAM_AWIDTH-1:0] bram_start_addr_for_inputs,
  input [`BRAM_AWIDTH-1:0] bram_start_addr_for_outputs
);

//addr mux
//one port on bram (a) is used by both external inputs and for writing results
//second port on bram (b) is used for reading inputs

wire [`BRAM_AWIDTH-1:0] bram_addr_a;
wire [`BRAM_AWIDTH-1:0] bram_addr_a_internal;
wire [`BRAM_AWIDTH-1:0] bram_addr_b;
wire [`BRAM_DWIDTH-1:0] bram_rdata_a;
wire [`BRAM_DWIDTH-1:0] bram_rdata_a_internal;
wire [`BRAM_DWIDTH-1:0] bram_rdata_b;
wire [`BRAM_DWIDTH-1:0] bram_wdata_a;
wire [`BRAM_DWIDTH-1:0] bram_wdata_a_internal;
wire [`BRAM_DWIDTH-1:0] bram_wdata_b;
wire bram_wren_a;
wire bram_wren_a_internal;
wire bram_wren_b;

wire [`NUM*`COMPUTE_DWIDTH-1:0] inp;
wire [31:0] out;

assign bram_wren_a = external ? bram_wren_ext : bram_wren_a_internal;
assign bram_wdata_a = external ? bram_wdata_ext : bram_wdata_a_internal;
assign bram_addr_a = external ? bram_addr_ext : bram_addr_a_internal;
assign bram_rdata_ext = bram_rdata_a;
assign bram_rdata_a_internal = bram_rdata_a;

assign bram_wren_b = ~bram_wren_a_internal;
assign bram_wdata_b = 0;

//instantiate bram
dpram u_ram(
    .clk(clk),
    .address_a(bram_addr_a),
    .address_b(bram_addr_b),
    .wren_a(bram_wren_a),
    .wren_b(bram_wren_b),
    .data_a(bram_wdata_a),
    .data_b(bram_wdata_b),
    .out_a(bram_rdata_a),
    .out_b(bram_rdata_b)
    );

//instantiate control logic
control_logic u_ctrl(
  .clk(clk),
  .reset(reset),
  .start(start),
  .done(done),
  .bram_start_addr_for_inputs(bram_start_addr_for_inputs),
  .bram_addr_for_inputs(bram_addr_b),
  .bram_data_inputs(bram_rdata_b),
  .bram_start_addr_for_outputs(bram_start_addr_for_outputs),
  .bram_addr_for_outputs(bram_addr_a_internal),
  .bram_data_outputs(bram_wdata_a_internal),
  .bram_we(bram_wren_a_internal),
  .inp(inp),
  .out(out)
);

//instantiate cu
compute_unit u_cu(
    .clk(clk),
    .reset(reset),
    .inp(inp),
    .out(out)
);

endmodule



module dpram (	
input clk,
input [`BRAM_AWIDTH-1:0] address_a,
input [`BRAM_AWIDTH-1:0] address_b,
input  wren_a,
input  wren_b,
input [`BRAM_DWIDTH-1:0] data_a,
input [`BRAM_DWIDTH-1:0] data_b,
output reg [`BRAM_DWIDTH-1:0] out_a,
output reg [`BRAM_DWIDTH-1:0] out_b
);


`ifdef VCS 

reg [`BRAM_DWIDTH-1:0] ram[`BRAM_DEPTH-1:0];

always @ (posedge clk) begin 
  if (wren_a) begin
      ram[address_a] <= data_a;
  end
  else begin
      out_a <= ram[address_a];
  end
end
  
always @ (posedge clk) begin 
  if (wren_b) begin
      ram[address_b] <= data_b;
  end 
  else begin
      out_b <= ram[address_b];
  end
end

`else

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif

`ifdef VCS
initial begin
  $vcdpluson;
  $vcdplusmemon;
end
`endif

endmodule



`define COMPUTE_DWIDTH 4
`define NUM 10
module compute_unit(
  input clk,
  input reset,
  input [`NUM*`COMPUTE_DWIDTH-1:0] inp,
  output [31:0] out
);

reg [`NUM*`COMPUTE_DWIDTH-1:0] input_reg;

always @(posedge clk) begin
    if (reset) begin
        input_reg <= 0;
    end 
    else begin
        input_reg <= inp;
    end    
end

wire [7:0] prod0;
wire [7:0] prod1;
wire [7:0] prod2;
wire [7:0] prod3;
wire [7:0] prod4;

assign prod0 = input_reg[7:4]   * input_reg[3:0];
assign prod1 = input_reg[15:12] * input_reg[11:8];
assign prod2 = input_reg[23:20] * input_reg[19:16];
assign prod3 = input_reg[31:28] * input_reg[27:24];
assign prod4 = input_reg[39:36] * input_reg[35:32];

reg [7:0] prod0_reg;
reg [7:0] prod1_reg;
reg [7:0] prod2_reg;
reg [7:0] prod3_reg;
reg [7:0] prod4_reg;

always @(posedge clk) begin
    if (reset) begin
        prod0_reg <= 0;
        prod1_reg <= 0;
        prod2_reg <= 0;
        prod3_reg <= 0;
        prod4_reg <= 0;
    end 
    else begin
        prod0_reg <= prod0;
        prod1_reg <= prod1;
        prod2_reg <= prod2;
        prod3_reg <= prod3;
        prod4_reg <= prod4;
    end    
end

wire [31:0] add1;
wire [31:0] add2;

assign add1 = prod0_reg + prod1_reg;
assign add2 = prod2_reg + prod3_reg;

reg [31:0] add1_reg;
reg [31:0] add2_reg;
reg [7:0] prod4_temp_reg;

always @(posedge clk) begin
    if (reset) begin
        add1_reg <= 0;
        add2_reg <= 0;
        prod4_temp_reg <= 0;
    end 
    else begin
        add1_reg <= add1;
        add2_reg <= add2;
        prod4_temp_reg <= prod4_reg;
    end    
end

wire [31:0] add3;

assign add3 = add1_reg + add2_reg;

reg [31:0] add3_reg;
reg [7:0] prod4_temp2_reg;

always @(posedge clk) begin
    if (reset) begin
        add3_reg <= 0;
        prod4_temp2_reg <= 0;
    end 
    else begin
        add3_reg <= add3;
        prod4_temp2_reg <= prod4_temp_reg;
    end    
end

wire [31:0] add4;

assign add4 = add3_reg + prod4_temp2_reg;

reg [31:0] add4_reg;

always @(posedge clk) begin
    if (reset) begin
        add4_reg <= 0;
    end 
    else begin
        add4_reg <= add4;
    end    
end

assign out = add4_reg;

endmodule

`define BRAM_DWIDTH 40
`define BRAM_AWIDTH 9
`define COMPUTE_DWIDTH 4
`define NUM 10

module control_logic(
  input clk,
  input reset,
  input start,
  output reg done,
  
  //bram interface
  input  [`BRAM_AWIDTH-1:0] bram_start_addr_for_inputs,
  output reg [`BRAM_AWIDTH-1:0] bram_addr_for_inputs,
  input  [`BRAM_DWIDTH-1:0] bram_data_inputs,
  input  [`BRAM_AWIDTH-1:0] bram_start_addr_for_outputs,
  output [`BRAM_AWIDTH-1:0] bram_addr_for_outputs,
  output [`BRAM_DWIDTH-1:0] bram_data_outputs,
  output reg bram_we,
  
  //interface with dot product unit
  output [`NUM*`COMPUTE_DWIDTH-1:0] inp,
  input  [31:0] out
);

reg [7:0] clk_cnt;
wire [9:0] clk_cnt_for_done;
assign clk_cnt_for_done = 472;

always @(posedge clk) begin
  if (reset || ~start) begin
    clk_cnt <= 0;
    done <= 0;
  end
  else if (clk_cnt == clk_cnt_for_done) begin
    done <= 1;
    clk_cnt <= clk_cnt + 1;
  end
  else if (done == 0) begin
    clk_cnt <= clk_cnt + 1;
  end    
  else begin
    done <= 0;
    clk_cnt <= clk_cnt + 1;
  end
end

//Reading inputs from BRAM
always @(posedge clk) begin
  if ((reset || ~start)) begin
    bram_addr_for_inputs <= bram_start_addr_for_inputs;
  end
  else begin
    bram_addr_for_inputs <= bram_addr_for_inputs + 1;
  end
end  

assign inp = bram_data_inputs;
assign bram_addr_for_outputs = bram_start_addr_for_outputs;

//Writing results to BRAM
always @(posedge clk) begin
  if ((reset || ~start || (clk_cnt == 472))) begin
    bram_we <= 1'b0;
  end
  else begin
    bram_we <= 1'b1;
  end
end  

assign bram_data_outputs = {8'b0,out};

endmodule
